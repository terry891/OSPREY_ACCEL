module CScratchpadPackedSubwordLoader(
  input          clock,
  input          reset,
  output         io_cache_block_in_ready,
  input          io_cache_block_in_valid,
  input  [511:0] io_cache_block_in_bits_dat,
  input  [6:0]   io_cache_block_in_bits_len,
  input  [5:0]   io_cache_block_in_bits_idxBase,
  output         io_sp_write_out_valid,
  output [127:0] io_sp_write_out_bits_dat,
  output [5:0]   io_sp_write_out_bits_idx
);
  reg [511:0] beat; // @[CScratchpadPackedSubwordLoader.scala 16:17]
  reg [5:0] idxBase; // @[CScratchpadPackedSubwordLoader.scala 17:20]
  reg [6:0] lenRemainingFromReq; // @[CScratchpadPackedSubwordLoader.scala 18:32]
  reg  state; // @[CScratchpadPackedSubwordLoader.scala 21:22]
  wire  _io_cache_block_in_ready_T = ~state; // @[CScratchpadPackedSubwordLoader.scala 22:36]
  wire  _T_1 = io_cache_block_in_ready & io_cache_block_in_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_0 = _T_1 | state; // @[CScratchpadPackedSubwordLoader.scala 34:36 35:15 21:22]
  wire [5:0] _idxBase_T_1 = idxBase + 6'h1; // @[CScratchpadPackedSubwordLoader.scala 50:28]
  wire [6:0] _lenRemainingFromReq_T_1 = lenRemainingFromReq - 7'h10; // @[CScratchpadPackedSubwordLoader.scala 53:54]
  wire  _GEN_6 = lenRemainingFromReq == 7'h10 ? 1'h0 : state; // @[CScratchpadPackedSubwordLoader.scala 54:60 55:19 21:22]
  wire [511:0] _GEN_10 = {{128'd0}, beat[511:128]}; // @[CScratchpadPackedSubwordLoader.scala 51:59 57:16 16:17]
  assign io_cache_block_in_ready = ~state; // @[CScratchpadPackedSubwordLoader.scala 22:36]
  assign io_sp_write_out_valid = _io_cache_block_in_ready_T ? 1'h0 : state; // @[CScratchpadPackedSubwordLoader.scala 32:17 24:25]
  assign io_sp_write_out_bits_dat = beat[127:0]; // @[CScratchpadPackedSubwordLoader.scala 29:9]
  assign io_sp_write_out_bits_idx = idxBase; // @[CScratchpadPackedSubwordLoader.scala 32:17 47:32]
  always @(posedge clock) begin
    if (_io_cache_block_in_ready_T) begin // @[CScratchpadPackedSubwordLoader.scala 32:17]
      if (_T_1) begin // @[CScratchpadPackedSubwordLoader.scala 34:36]
        beat <= io_cache_block_in_bits_dat; // @[CScratchpadPackedSubwordLoader.scala 36:14]
      end
    end else if (state) begin // @[CScratchpadPackedSubwordLoader.scala 32:17]
      if (io_sp_write_out_valid) begin // @[CScratchpadPackedSubwordLoader.scala 48:34]
        beat <= _GEN_10;
      end
    end
    if (_io_cache_block_in_ready_T) begin // @[CScratchpadPackedSubwordLoader.scala 32:17]
      if (_T_1) begin // @[CScratchpadPackedSubwordLoader.scala 34:36]
        idxBase <= io_cache_block_in_bits_idxBase; // @[CScratchpadPackedSubwordLoader.scala 37:17]
      end
    end else if (state) begin // @[CScratchpadPackedSubwordLoader.scala 32:17]
      if (io_sp_write_out_valid) begin // @[CScratchpadPackedSubwordLoader.scala 48:34]
        idxBase <= _idxBase_T_1; // @[CScratchpadPackedSubwordLoader.scala 50:17]
      end
    end
    if (_io_cache_block_in_ready_T) begin // @[CScratchpadPackedSubwordLoader.scala 32:17]
      if (_T_1) begin // @[CScratchpadPackedSubwordLoader.scala 34:36]
        lenRemainingFromReq <= io_cache_block_in_bits_len; // @[CScratchpadPackedSubwordLoader.scala 38:29]
      end
    end else if (state) begin // @[CScratchpadPackedSubwordLoader.scala 32:17]
      if (io_sp_write_out_valid) begin // @[CScratchpadPackedSubwordLoader.scala 48:34]
        lenRemainingFromReq <= _lenRemainingFromReq_T_1;
      end
    end
    if (reset) begin // @[CScratchpadPackedSubwordLoader.scala 21:22]
      state <= 1'h0; // @[CScratchpadPackedSubwordLoader.scala 21:22]
    end else if (_io_cache_block_in_ready_T) begin // @[CScratchpadPackedSubwordLoader.scala 32:17]
      state <= _GEN_0;
    end else if (state) begin // @[CScratchpadPackedSubwordLoader.scala 32:17]
      if (io_sp_write_out_valid) begin // @[CScratchpadPackedSubwordLoader.scala 48:34]
        state <= _GEN_6;
      end
    end
  end
endmodule
module CScratchpad(
  input          clock,
  input          reset,
  input          auto_mem_out_a_ready,
  output         auto_mem_out_a_valid,
  output [2:0]   auto_mem_out_a_bits_size,
  output [3:0]   auto_mem_out_a_bits_source,
  output [33:0]  auto_mem_out_a_bits_address,
  output [63:0]  auto_mem_out_a_bits_mask,
  output         auto_mem_out_d_ready,
  input          auto_mem_out_d_valid,
  input  [3:0]   auto_mem_out_d_bits_source,
  input  [511:0] auto_mem_out_d_bits_data,
  input          access_readReq_valid,
  output         access_readRes_valid,
  output [127:0] access_readRes_bits
);
  reg [127:0] mem [0:63]; // @[CScratchpad.scala 92:24]
  wire  mem_rval_en; // @[CScratchpad.scala 92:24]
  wire [5:0] mem_rval_addr; // @[CScratchpad.scala 92:24]
  wire [127:0] mem_rval_data; // @[CScratchpad.scala 92:24]
  wire [127:0] mem_MPORT_data; // @[CScratchpad.scala 92:24]
  wire [5:0] mem_MPORT_addr; // @[CScratchpad.scala 92:24]
  wire  mem_MPORT_mask; // @[CScratchpad.scala 92:24]
  wire  mem_MPORT_en; // @[CScratchpad.scala 92:24]
  wire [127:0] mem_MPORT_1_data; // @[CScratchpad.scala 92:24]
  wire [5:0] mem_MPORT_1_addr; // @[CScratchpad.scala 92:24]
  wire  mem_MPORT_1_mask; // @[CScratchpad.scala 92:24]
  wire  mem_MPORT_1_en; // @[CScratchpad.scala 92:24]
  reg  mem_rval_en_pipe_0;
  reg [5:0] mem_rval_addr_pipe_0;
  wire  loader_clock; // @[CScratchpad.scala 94:30]
  wire  loader_reset; // @[CScratchpad.scala 94:30]
  wire  loader_io_cache_block_in_ready; // @[CScratchpad.scala 94:30]
  wire  loader_io_cache_block_in_valid; // @[CScratchpad.scala 94:30]
  wire [511:0] loader_io_cache_block_in_bits_dat; // @[CScratchpad.scala 94:30]
  wire [6:0] loader_io_cache_block_in_bits_len; // @[CScratchpad.scala 94:30]
  wire [5:0] loader_io_cache_block_in_bits_idxBase; // @[CScratchpad.scala 94:30]
  wire  loader_io_sp_write_out_valid; // @[CScratchpad.scala 94:30]
  wire [127:0] loader_io_sp_write_out_bits_dat; // @[CScratchpad.scala 94:30]
  wire [5:0] loader_io_sp_write_out_bits_idx; // @[CScratchpad.scala 94:30]
  reg [1:0] mem_tx_state; // @[CScratchpad.scala 102:37]
  reg  access_readRes_valid_REG; // @[CScratchpad.scala 85:30]
  reg  reqIdleBits_0; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_1; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_2; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_3; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_4; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_5; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_6; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_7; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_8; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_9; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_10; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_11; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_12; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_13; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_14; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_15; // @[CScratchpad.scala 110:36]
  wire  reqAvailable = reqIdleBits_0 | reqIdleBits_1 | reqIdleBits_2 | reqIdleBits_3 | reqIdleBits_4 | reqIdleBits_5 |
    reqIdleBits_6 | reqIdleBits_7 | reqIdleBits_8 | reqIdleBits_9 | reqIdleBits_10 | reqIdleBits_11 | reqIdleBits_12 |
    reqIdleBits_13 | reqIdleBits_14 | reqIdleBits_15; // @[CScratchpad.scala 111:51]
  wire [3:0] _reqChosen_T = reqIdleBits_14 ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_1 = reqIdleBits_13 ? 4'hd : _reqChosen_T; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_2 = reqIdleBits_12 ? 4'hc : _reqChosen_T_1; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_3 = reqIdleBits_11 ? 4'hb : _reqChosen_T_2; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_4 = reqIdleBits_10 ? 4'ha : _reqChosen_T_3; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_5 = reqIdleBits_9 ? 4'h9 : _reqChosen_T_4; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_6 = reqIdleBits_8 ? 4'h8 : _reqChosen_T_5; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_7 = reqIdleBits_7 ? 4'h7 : _reqChosen_T_6; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_8 = reqIdleBits_6 ? 4'h6 : _reqChosen_T_7; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_9 = reqIdleBits_5 ? 4'h5 : _reqChosen_T_8; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_10 = reqIdleBits_4 ? 4'h4 : _reqChosen_T_9; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_11 = reqIdleBits_3 ? 4'h3 : _reqChosen_T_10; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_12 = reqIdleBits_2 ? 4'h2 : _reqChosen_T_11; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_13 = reqIdleBits_1 ? 4'h1 : _reqChosen_T_12; // @[Mux.scala 47:70]
  wire [3:0] reqChosen = reqIdleBits_0 ? 4'h0 : _reqChosen_T_13; // @[Mux.scala 47:70]
  reg [5:0] req_cache_0_scratchpadAddress; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_0_memoryLength; // @[CScratchpad.scala 114:30]
  reg [5:0] req_cache_1_scratchpadAddress; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_1_memoryLength; // @[CScratchpad.scala 114:30]
  reg [5:0] req_cache_2_scratchpadAddress; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_2_memoryLength; // @[CScratchpad.scala 114:30]
  reg [5:0] req_cache_3_scratchpadAddress; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_3_memoryLength; // @[CScratchpad.scala 114:30]
  reg [5:0] req_cache_4_scratchpadAddress; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_4_memoryLength; // @[CScratchpad.scala 114:30]
  reg [5:0] req_cache_5_scratchpadAddress; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_5_memoryLength; // @[CScratchpad.scala 114:30]
  reg [5:0] req_cache_6_scratchpadAddress; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_6_memoryLength; // @[CScratchpad.scala 114:30]
  reg [5:0] req_cache_7_scratchpadAddress; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_7_memoryLength; // @[CScratchpad.scala 114:30]
  reg [5:0] req_cache_8_scratchpadAddress; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_8_memoryLength; // @[CScratchpad.scala 114:30]
  reg [5:0] req_cache_9_scratchpadAddress; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_9_memoryLength; // @[CScratchpad.scala 114:30]
  reg [5:0] req_cache_10_scratchpadAddress; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_10_memoryLength; // @[CScratchpad.scala 114:30]
  reg [5:0] req_cache_11_scratchpadAddress; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_11_memoryLength; // @[CScratchpad.scala 114:30]
  reg [5:0] req_cache_12_scratchpadAddress; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_12_memoryLength; // @[CScratchpad.scala 114:30]
  reg [5:0] req_cache_13_scratchpadAddress; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_13_memoryLength; // @[CScratchpad.scala 114:30]
  reg [5:0] req_cache_14_scratchpadAddress; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_14_memoryLength; // @[CScratchpad.scala 114:30]
  reg [5:0] req_cache_15_scratchpadAddress; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_15_memoryLength; // @[CScratchpad.scala 114:30]
  reg [33:0] totalTx_memoryAddress; // @[CScratchpad.scala 124:28]
  reg [5:0] totalTx_scratchpadAddress; // @[CScratchpad.scala 124:28]
  reg [33:0] totalTx_memoryLength; // @[CScratchpad.scala 124:28]
  wire  isBelowLimit = totalTx_memoryLength <= 34'h40; // @[CScratchpad.scala 149:47]
  wire [1:0] txEmitLengthLg_hi = totalTx_memoryLength[33:32]; // @[OneHot.scala 30:18]
  wire  _txEmitLengthLg_T = |txEmitLengthLg_hi; // @[OneHot.scala 32:14]
  wire [31:0] txEmitLengthLg_lo = totalTx_memoryLength[31:0]; // @[OneHot.scala 31:18]
  wire [31:0] _GEN_569 = {{30'd0}, txEmitLengthLg_hi}; // @[OneHot.scala 32:28]
  wire [31:0] _txEmitLengthLg_T_1 = _GEN_569 | txEmitLengthLg_lo; // @[OneHot.scala 32:28]
  wire [15:0] txEmitLengthLg_hi_1 = _txEmitLengthLg_T_1[31:16]; // @[OneHot.scala 30:18]
  wire  _txEmitLengthLg_T_2 = |txEmitLengthLg_hi_1; // @[OneHot.scala 32:14]
  wire [15:0] txEmitLengthLg_lo_1 = _txEmitLengthLg_T_1[15:0]; // @[OneHot.scala 31:18]
  wire [15:0] _txEmitLengthLg_T_3 = txEmitLengthLg_hi_1 | txEmitLengthLg_lo_1; // @[OneHot.scala 32:28]
  wire [7:0] txEmitLengthLg_hi_2 = _txEmitLengthLg_T_3[15:8]; // @[OneHot.scala 30:18]
  wire  _txEmitLengthLg_T_4 = |txEmitLengthLg_hi_2; // @[OneHot.scala 32:14]
  wire [7:0] txEmitLengthLg_lo_2 = _txEmitLengthLg_T_3[7:0]; // @[OneHot.scala 31:18]
  wire [7:0] _txEmitLengthLg_T_5 = txEmitLengthLg_hi_2 | txEmitLengthLg_lo_2; // @[OneHot.scala 32:28]
  wire [3:0] txEmitLengthLg_hi_3 = _txEmitLengthLg_T_5[7:4]; // @[OneHot.scala 30:18]
  wire  _txEmitLengthLg_T_6 = |txEmitLengthLg_hi_3; // @[OneHot.scala 32:14]
  wire [3:0] txEmitLengthLg_lo_3 = _txEmitLengthLg_T_5[3:0]; // @[OneHot.scala 31:18]
  wire [3:0] _txEmitLengthLg_T_7 = txEmitLengthLg_hi_3 | txEmitLengthLg_lo_3; // @[OneHot.scala 32:28]
  wire [1:0] txEmitLengthLg_hi_4 = _txEmitLengthLg_T_7[3:2]; // @[OneHot.scala 30:18]
  wire  _txEmitLengthLg_T_8 = |txEmitLengthLg_hi_4; // @[OneHot.scala 32:14]
  wire [1:0] txEmitLengthLg_lo_4 = _txEmitLengthLg_T_7[1:0]; // @[OneHot.scala 31:18]
  wire [1:0] _txEmitLengthLg_T_9 = txEmitLengthLg_hi_4 | txEmitLengthLg_lo_4; // @[OneHot.scala 32:28]
  wire [5:0] _txEmitLengthLg_T_15 = {_txEmitLengthLg_T,_txEmitLengthLg_T_2,_txEmitLengthLg_T_4,_txEmitLengthLg_T_6,
    _txEmitLengthLg_T_8,_txEmitLengthLg_T_9[1]}; // @[Cat.scala 33:92]
  wire [5:0] _txEmitLengthLg_T_16 = isBelowLimit ? _txEmitLengthLg_T_15 : 6'h6; // @[CScratchpad.scala 150:28]
  wire [5:0] _GEN_111 = 2'h1 == mem_tx_state ? _txEmitLengthLg_T_16 : 6'h0; // @[CScratchpad.scala 131:18 138:24 150:22]
  wire [5:0] _GEN_169 = 2'h0 == mem_tx_state ? 6'h0 : _GEN_111; // @[CScratchpad.scala 131:18 138:24]
  wire [3:0] txEmitLengthLg = _GEN_169[3:0]; // @[CScratchpad.scala 130:36]
  wire [5:0] _x1_a_bits_a_mask_sizeOH_T = {{2'd0}, txEmitLengthLg}; // @[Misc.scala 201:34]
  wire [2:0] x1_a_bits_a_mask_sizeOH_shiftAmount = _x1_a_bits_a_mask_sizeOH_T[2:0]; // @[OneHot.scala 63:49]
  wire [7:0] _x1_a_bits_a_mask_sizeOH_T_1 = 8'h1 << x1_a_bits_a_mask_sizeOH_shiftAmount; // @[OneHot.scala 64:12]
  wire [5:0] x1_a_bits_a_mask_sizeOH = _x1_a_bits_a_mask_sizeOH_T_1[5:0] | 6'h1; // @[Misc.scala 201:81]
  wire  _x1_a_bits_a_mask_T = txEmitLengthLg >= 4'h6; // @[Misc.scala 205:21]
  wire  x1_a_bits_a_mask_size = x1_a_bits_a_mask_sizeOH[5]; // @[Misc.scala 208:26]
  wire  x1_a_bits_a_mask_bit = totalTx_memoryAddress[5]; // @[Misc.scala 209:26]
  wire  x1_a_bits_a_mask_nbit = ~x1_a_bits_a_mask_bit; // @[Misc.scala 210:20]
  wire  x1_a_bits_a_mask_acc = _x1_a_bits_a_mask_T | x1_a_bits_a_mask_size & x1_a_bits_a_mask_nbit; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_acc_1 = _x1_a_bits_a_mask_T | x1_a_bits_a_mask_size & x1_a_bits_a_mask_bit; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_size_1 = x1_a_bits_a_mask_sizeOH[4]; // @[Misc.scala 208:26]
  wire  x1_a_bits_a_mask_bit_1 = totalTx_memoryAddress[4]; // @[Misc.scala 209:26]
  wire  x1_a_bits_a_mask_nbit_1 = ~x1_a_bits_a_mask_bit_1; // @[Misc.scala 210:20]
  wire  x1_a_bits_a_mask_eq_2 = x1_a_bits_a_mask_nbit & x1_a_bits_a_mask_nbit_1; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_2 = x1_a_bits_a_mask_acc | x1_a_bits_a_mask_size_1 & x1_a_bits_a_mask_eq_2; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_3 = x1_a_bits_a_mask_nbit & x1_a_bits_a_mask_bit_1; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_3 = x1_a_bits_a_mask_acc | x1_a_bits_a_mask_size_1 & x1_a_bits_a_mask_eq_3; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_4 = x1_a_bits_a_mask_bit & x1_a_bits_a_mask_nbit_1; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_4 = x1_a_bits_a_mask_acc_1 | x1_a_bits_a_mask_size_1 & x1_a_bits_a_mask_eq_4; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_5 = x1_a_bits_a_mask_bit & x1_a_bits_a_mask_bit_1; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_5 = x1_a_bits_a_mask_acc_1 | x1_a_bits_a_mask_size_1 & x1_a_bits_a_mask_eq_5; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_size_2 = x1_a_bits_a_mask_sizeOH[3]; // @[Misc.scala 208:26]
  wire  x1_a_bits_a_mask_bit_2 = totalTx_memoryAddress[3]; // @[Misc.scala 209:26]
  wire  x1_a_bits_a_mask_nbit_2 = ~x1_a_bits_a_mask_bit_2; // @[Misc.scala 210:20]
  wire  x1_a_bits_a_mask_eq_6 = x1_a_bits_a_mask_eq_2 & x1_a_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_6 = x1_a_bits_a_mask_acc_2 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_6; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_7 = x1_a_bits_a_mask_eq_2 & x1_a_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_7 = x1_a_bits_a_mask_acc_2 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_7; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_8 = x1_a_bits_a_mask_eq_3 & x1_a_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_8 = x1_a_bits_a_mask_acc_3 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_8; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_9 = x1_a_bits_a_mask_eq_3 & x1_a_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_9 = x1_a_bits_a_mask_acc_3 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_9; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_10 = x1_a_bits_a_mask_eq_4 & x1_a_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_10 = x1_a_bits_a_mask_acc_4 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_10; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_11 = x1_a_bits_a_mask_eq_4 & x1_a_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_11 = x1_a_bits_a_mask_acc_4 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_11; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_12 = x1_a_bits_a_mask_eq_5 & x1_a_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_12 = x1_a_bits_a_mask_acc_5 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_12; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_13 = x1_a_bits_a_mask_eq_5 & x1_a_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_13 = x1_a_bits_a_mask_acc_5 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_13; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_size_3 = x1_a_bits_a_mask_sizeOH[2]; // @[Misc.scala 208:26]
  wire  x1_a_bits_a_mask_bit_3 = totalTx_memoryAddress[2]; // @[Misc.scala 209:26]
  wire  x1_a_bits_a_mask_nbit_3 = ~x1_a_bits_a_mask_bit_3; // @[Misc.scala 210:20]
  wire  x1_a_bits_a_mask_eq_14 = x1_a_bits_a_mask_eq_6 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_14 = x1_a_bits_a_mask_acc_6 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_14; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_15 = x1_a_bits_a_mask_eq_6 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_15 = x1_a_bits_a_mask_acc_6 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_15; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_16 = x1_a_bits_a_mask_eq_7 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_16 = x1_a_bits_a_mask_acc_7 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_16; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_17 = x1_a_bits_a_mask_eq_7 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_17 = x1_a_bits_a_mask_acc_7 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_17; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_18 = x1_a_bits_a_mask_eq_8 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_18 = x1_a_bits_a_mask_acc_8 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_18; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_19 = x1_a_bits_a_mask_eq_8 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_19 = x1_a_bits_a_mask_acc_8 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_19; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_20 = x1_a_bits_a_mask_eq_9 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_20 = x1_a_bits_a_mask_acc_9 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_20; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_21 = x1_a_bits_a_mask_eq_9 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_21 = x1_a_bits_a_mask_acc_9 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_21; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_22 = x1_a_bits_a_mask_eq_10 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_22 = x1_a_bits_a_mask_acc_10 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_22; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_23 = x1_a_bits_a_mask_eq_10 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_23 = x1_a_bits_a_mask_acc_10 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_23; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_24 = x1_a_bits_a_mask_eq_11 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_24 = x1_a_bits_a_mask_acc_11 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_24; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_25 = x1_a_bits_a_mask_eq_11 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_25 = x1_a_bits_a_mask_acc_11 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_25; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_26 = x1_a_bits_a_mask_eq_12 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_26 = x1_a_bits_a_mask_acc_12 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_26; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_27 = x1_a_bits_a_mask_eq_12 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_27 = x1_a_bits_a_mask_acc_12 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_27; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_28 = x1_a_bits_a_mask_eq_13 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_28 = x1_a_bits_a_mask_acc_13 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_28; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_29 = x1_a_bits_a_mask_eq_13 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_29 = x1_a_bits_a_mask_acc_13 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_29; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_size_4 = x1_a_bits_a_mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  x1_a_bits_a_mask_bit_4 = totalTx_memoryAddress[1]; // @[Misc.scala 209:26]
  wire  x1_a_bits_a_mask_nbit_4 = ~x1_a_bits_a_mask_bit_4; // @[Misc.scala 210:20]
  wire  x1_a_bits_a_mask_eq_30 = x1_a_bits_a_mask_eq_14 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_30 = x1_a_bits_a_mask_acc_14 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_30; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_31 = x1_a_bits_a_mask_eq_14 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_31 = x1_a_bits_a_mask_acc_14 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_31; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_32 = x1_a_bits_a_mask_eq_15 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_32 = x1_a_bits_a_mask_acc_15 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_32; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_33 = x1_a_bits_a_mask_eq_15 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_33 = x1_a_bits_a_mask_acc_15 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_33; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_34 = x1_a_bits_a_mask_eq_16 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_34 = x1_a_bits_a_mask_acc_16 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_34; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_35 = x1_a_bits_a_mask_eq_16 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_35 = x1_a_bits_a_mask_acc_16 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_35; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_36 = x1_a_bits_a_mask_eq_17 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_36 = x1_a_bits_a_mask_acc_17 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_36; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_37 = x1_a_bits_a_mask_eq_17 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_37 = x1_a_bits_a_mask_acc_17 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_37; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_38 = x1_a_bits_a_mask_eq_18 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_38 = x1_a_bits_a_mask_acc_18 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_38; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_39 = x1_a_bits_a_mask_eq_18 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_39 = x1_a_bits_a_mask_acc_18 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_39; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_40 = x1_a_bits_a_mask_eq_19 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_40 = x1_a_bits_a_mask_acc_19 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_40; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_41 = x1_a_bits_a_mask_eq_19 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_41 = x1_a_bits_a_mask_acc_19 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_41; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_42 = x1_a_bits_a_mask_eq_20 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_42 = x1_a_bits_a_mask_acc_20 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_42; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_43 = x1_a_bits_a_mask_eq_20 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_43 = x1_a_bits_a_mask_acc_20 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_43; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_44 = x1_a_bits_a_mask_eq_21 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_44 = x1_a_bits_a_mask_acc_21 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_44; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_45 = x1_a_bits_a_mask_eq_21 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_45 = x1_a_bits_a_mask_acc_21 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_45; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_46 = x1_a_bits_a_mask_eq_22 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_46 = x1_a_bits_a_mask_acc_22 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_46; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_47 = x1_a_bits_a_mask_eq_22 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_47 = x1_a_bits_a_mask_acc_22 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_47; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_48 = x1_a_bits_a_mask_eq_23 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_48 = x1_a_bits_a_mask_acc_23 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_48; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_49 = x1_a_bits_a_mask_eq_23 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_49 = x1_a_bits_a_mask_acc_23 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_49; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_50 = x1_a_bits_a_mask_eq_24 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_50 = x1_a_bits_a_mask_acc_24 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_50; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_51 = x1_a_bits_a_mask_eq_24 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_51 = x1_a_bits_a_mask_acc_24 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_51; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_52 = x1_a_bits_a_mask_eq_25 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_52 = x1_a_bits_a_mask_acc_25 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_52; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_53 = x1_a_bits_a_mask_eq_25 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_53 = x1_a_bits_a_mask_acc_25 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_53; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_54 = x1_a_bits_a_mask_eq_26 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_54 = x1_a_bits_a_mask_acc_26 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_54; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_55 = x1_a_bits_a_mask_eq_26 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_55 = x1_a_bits_a_mask_acc_26 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_55; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_56 = x1_a_bits_a_mask_eq_27 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_56 = x1_a_bits_a_mask_acc_27 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_56; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_57 = x1_a_bits_a_mask_eq_27 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_57 = x1_a_bits_a_mask_acc_27 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_57; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_58 = x1_a_bits_a_mask_eq_28 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_58 = x1_a_bits_a_mask_acc_28 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_58; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_59 = x1_a_bits_a_mask_eq_28 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_59 = x1_a_bits_a_mask_acc_28 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_59; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_60 = x1_a_bits_a_mask_eq_29 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_60 = x1_a_bits_a_mask_acc_29 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_60; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_61 = x1_a_bits_a_mask_eq_29 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_61 = x1_a_bits_a_mask_acc_29 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_61; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_size_5 = x1_a_bits_a_mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  x1_a_bits_a_mask_bit_5 = totalTx_memoryAddress[0]; // @[Misc.scala 209:26]
  wire  x1_a_bits_a_mask_nbit_5 = ~x1_a_bits_a_mask_bit_5; // @[Misc.scala 210:20]
  wire  x1_a_bits_a_mask_eq_62 = x1_a_bits_a_mask_eq_30 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_62 = x1_a_bits_a_mask_acc_30 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_62; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_63 = x1_a_bits_a_mask_eq_30 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_63 = x1_a_bits_a_mask_acc_30 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_63; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_64 = x1_a_bits_a_mask_eq_31 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_64 = x1_a_bits_a_mask_acc_31 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_64; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_65 = x1_a_bits_a_mask_eq_31 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_65 = x1_a_bits_a_mask_acc_31 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_65; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_66 = x1_a_bits_a_mask_eq_32 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_66 = x1_a_bits_a_mask_acc_32 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_66; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_67 = x1_a_bits_a_mask_eq_32 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_67 = x1_a_bits_a_mask_acc_32 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_67; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_68 = x1_a_bits_a_mask_eq_33 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_68 = x1_a_bits_a_mask_acc_33 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_68; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_69 = x1_a_bits_a_mask_eq_33 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_69 = x1_a_bits_a_mask_acc_33 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_69; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_70 = x1_a_bits_a_mask_eq_34 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_70 = x1_a_bits_a_mask_acc_34 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_70; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_71 = x1_a_bits_a_mask_eq_34 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_71 = x1_a_bits_a_mask_acc_34 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_71; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_72 = x1_a_bits_a_mask_eq_35 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_72 = x1_a_bits_a_mask_acc_35 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_72; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_73 = x1_a_bits_a_mask_eq_35 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_73 = x1_a_bits_a_mask_acc_35 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_73; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_74 = x1_a_bits_a_mask_eq_36 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_74 = x1_a_bits_a_mask_acc_36 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_74; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_75 = x1_a_bits_a_mask_eq_36 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_75 = x1_a_bits_a_mask_acc_36 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_75; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_76 = x1_a_bits_a_mask_eq_37 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_76 = x1_a_bits_a_mask_acc_37 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_76; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_77 = x1_a_bits_a_mask_eq_37 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_77 = x1_a_bits_a_mask_acc_37 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_77; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_78 = x1_a_bits_a_mask_eq_38 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_78 = x1_a_bits_a_mask_acc_38 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_78; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_79 = x1_a_bits_a_mask_eq_38 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_79 = x1_a_bits_a_mask_acc_38 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_79; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_80 = x1_a_bits_a_mask_eq_39 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_80 = x1_a_bits_a_mask_acc_39 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_80; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_81 = x1_a_bits_a_mask_eq_39 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_81 = x1_a_bits_a_mask_acc_39 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_81; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_82 = x1_a_bits_a_mask_eq_40 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_82 = x1_a_bits_a_mask_acc_40 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_82; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_83 = x1_a_bits_a_mask_eq_40 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_83 = x1_a_bits_a_mask_acc_40 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_83; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_84 = x1_a_bits_a_mask_eq_41 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_84 = x1_a_bits_a_mask_acc_41 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_84; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_85 = x1_a_bits_a_mask_eq_41 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_85 = x1_a_bits_a_mask_acc_41 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_85; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_86 = x1_a_bits_a_mask_eq_42 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_86 = x1_a_bits_a_mask_acc_42 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_86; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_87 = x1_a_bits_a_mask_eq_42 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_87 = x1_a_bits_a_mask_acc_42 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_87; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_88 = x1_a_bits_a_mask_eq_43 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_88 = x1_a_bits_a_mask_acc_43 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_88; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_89 = x1_a_bits_a_mask_eq_43 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_89 = x1_a_bits_a_mask_acc_43 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_89; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_90 = x1_a_bits_a_mask_eq_44 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_90 = x1_a_bits_a_mask_acc_44 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_90; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_91 = x1_a_bits_a_mask_eq_44 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_91 = x1_a_bits_a_mask_acc_44 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_91; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_92 = x1_a_bits_a_mask_eq_45 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_92 = x1_a_bits_a_mask_acc_45 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_92; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_93 = x1_a_bits_a_mask_eq_45 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_93 = x1_a_bits_a_mask_acc_45 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_93; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_94 = x1_a_bits_a_mask_eq_46 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_94 = x1_a_bits_a_mask_acc_46 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_94; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_95 = x1_a_bits_a_mask_eq_46 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_95 = x1_a_bits_a_mask_acc_46 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_95; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_96 = x1_a_bits_a_mask_eq_47 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_96 = x1_a_bits_a_mask_acc_47 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_96; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_97 = x1_a_bits_a_mask_eq_47 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_97 = x1_a_bits_a_mask_acc_47 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_97; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_98 = x1_a_bits_a_mask_eq_48 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_98 = x1_a_bits_a_mask_acc_48 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_98; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_99 = x1_a_bits_a_mask_eq_48 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_99 = x1_a_bits_a_mask_acc_48 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_99; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_100 = x1_a_bits_a_mask_eq_49 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_100 = x1_a_bits_a_mask_acc_49 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_100; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_101 = x1_a_bits_a_mask_eq_49 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_101 = x1_a_bits_a_mask_acc_49 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_101; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_102 = x1_a_bits_a_mask_eq_50 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_102 = x1_a_bits_a_mask_acc_50 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_102; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_103 = x1_a_bits_a_mask_eq_50 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_103 = x1_a_bits_a_mask_acc_50 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_103; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_104 = x1_a_bits_a_mask_eq_51 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_104 = x1_a_bits_a_mask_acc_51 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_104; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_105 = x1_a_bits_a_mask_eq_51 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_105 = x1_a_bits_a_mask_acc_51 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_105; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_106 = x1_a_bits_a_mask_eq_52 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_106 = x1_a_bits_a_mask_acc_52 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_106; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_107 = x1_a_bits_a_mask_eq_52 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_107 = x1_a_bits_a_mask_acc_52 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_107; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_108 = x1_a_bits_a_mask_eq_53 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_108 = x1_a_bits_a_mask_acc_53 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_108; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_109 = x1_a_bits_a_mask_eq_53 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_109 = x1_a_bits_a_mask_acc_53 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_109; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_110 = x1_a_bits_a_mask_eq_54 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_110 = x1_a_bits_a_mask_acc_54 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_110; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_111 = x1_a_bits_a_mask_eq_54 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_111 = x1_a_bits_a_mask_acc_54 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_111; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_112 = x1_a_bits_a_mask_eq_55 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_112 = x1_a_bits_a_mask_acc_55 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_112; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_113 = x1_a_bits_a_mask_eq_55 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_113 = x1_a_bits_a_mask_acc_55 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_113; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_114 = x1_a_bits_a_mask_eq_56 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_114 = x1_a_bits_a_mask_acc_56 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_114; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_115 = x1_a_bits_a_mask_eq_56 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_115 = x1_a_bits_a_mask_acc_56 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_115; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_116 = x1_a_bits_a_mask_eq_57 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_116 = x1_a_bits_a_mask_acc_57 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_116; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_117 = x1_a_bits_a_mask_eq_57 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_117 = x1_a_bits_a_mask_acc_57 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_117; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_118 = x1_a_bits_a_mask_eq_58 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_118 = x1_a_bits_a_mask_acc_58 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_118; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_119 = x1_a_bits_a_mask_eq_58 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_119 = x1_a_bits_a_mask_acc_58 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_119; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_120 = x1_a_bits_a_mask_eq_59 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_120 = x1_a_bits_a_mask_acc_59 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_120; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_121 = x1_a_bits_a_mask_eq_59 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_121 = x1_a_bits_a_mask_acc_59 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_121; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_122 = x1_a_bits_a_mask_eq_60 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_122 = x1_a_bits_a_mask_acc_60 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_122; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_123 = x1_a_bits_a_mask_eq_60 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_123 = x1_a_bits_a_mask_acc_60 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_123; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_124 = x1_a_bits_a_mask_eq_61 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_124 = x1_a_bits_a_mask_acc_61 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_124; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_125 = x1_a_bits_a_mask_eq_61 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_125 = x1_a_bits_a_mask_acc_61 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_125; // @[Misc.scala 214:29]
  wire [7:0] x1_a_bits_a_mask_lo_lo_lo = {x1_a_bits_a_mask_acc_69,x1_a_bits_a_mask_acc_68,x1_a_bits_a_mask_acc_67,
    x1_a_bits_a_mask_acc_66,x1_a_bits_a_mask_acc_65,x1_a_bits_a_mask_acc_64,x1_a_bits_a_mask_acc_63,
    x1_a_bits_a_mask_acc_62}; // @[Cat.scala 33:92]
  wire [15:0] x1_a_bits_a_mask_lo_lo = {x1_a_bits_a_mask_acc_77,x1_a_bits_a_mask_acc_76,x1_a_bits_a_mask_acc_75,
    x1_a_bits_a_mask_acc_74,x1_a_bits_a_mask_acc_73,x1_a_bits_a_mask_acc_72,x1_a_bits_a_mask_acc_71,
    x1_a_bits_a_mask_acc_70,x1_a_bits_a_mask_lo_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] x1_a_bits_a_mask_lo_hi_lo = {x1_a_bits_a_mask_acc_85,x1_a_bits_a_mask_acc_84,x1_a_bits_a_mask_acc_83,
    x1_a_bits_a_mask_acc_82,x1_a_bits_a_mask_acc_81,x1_a_bits_a_mask_acc_80,x1_a_bits_a_mask_acc_79,
    x1_a_bits_a_mask_acc_78}; // @[Cat.scala 33:92]
  wire [31:0] x1_a_bits_a_mask_lo = {x1_a_bits_a_mask_acc_93,x1_a_bits_a_mask_acc_92,x1_a_bits_a_mask_acc_91,
    x1_a_bits_a_mask_acc_90,x1_a_bits_a_mask_acc_89,x1_a_bits_a_mask_acc_88,x1_a_bits_a_mask_acc_87,
    x1_a_bits_a_mask_acc_86,x1_a_bits_a_mask_lo_hi_lo,x1_a_bits_a_mask_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] x1_a_bits_a_mask_hi_lo_lo = {x1_a_bits_a_mask_acc_101,x1_a_bits_a_mask_acc_100,x1_a_bits_a_mask_acc_99,
    x1_a_bits_a_mask_acc_98,x1_a_bits_a_mask_acc_97,x1_a_bits_a_mask_acc_96,x1_a_bits_a_mask_acc_95,
    x1_a_bits_a_mask_acc_94}; // @[Cat.scala 33:92]
  wire [15:0] x1_a_bits_a_mask_hi_lo = {x1_a_bits_a_mask_acc_109,x1_a_bits_a_mask_acc_108,x1_a_bits_a_mask_acc_107,
    x1_a_bits_a_mask_acc_106,x1_a_bits_a_mask_acc_105,x1_a_bits_a_mask_acc_104,x1_a_bits_a_mask_acc_103,
    x1_a_bits_a_mask_acc_102,x1_a_bits_a_mask_hi_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] x1_a_bits_a_mask_hi_hi_lo = {x1_a_bits_a_mask_acc_117,x1_a_bits_a_mask_acc_116,x1_a_bits_a_mask_acc_115,
    x1_a_bits_a_mask_acc_114,x1_a_bits_a_mask_acc_113,x1_a_bits_a_mask_acc_112,x1_a_bits_a_mask_acc_111,
    x1_a_bits_a_mask_acc_110}; // @[Cat.scala 33:92]
  wire [31:0] x1_a_bits_a_mask_hi = {x1_a_bits_a_mask_acc_125,x1_a_bits_a_mask_acc_124,x1_a_bits_a_mask_acc_123,
    x1_a_bits_a_mask_acc_122,x1_a_bits_a_mask_acc_121,x1_a_bits_a_mask_acc_120,x1_a_bits_a_mask_acc_119,
    x1_a_bits_a_mask_acc_118,x1_a_bits_a_mask_hi_hi_lo,x1_a_bits_a_mask_hi_lo}; // @[Cat.scala 33:92]
  wire  _GEN_112 = 2'h1 == mem_tx_state ? reqAvailable : mem_tx_state == 2'h1; // @[CScratchpad.scala 136:19 138:24 151:23]
  wire  mem_out_a_valid = 2'h0 == mem_tx_state ? mem_tx_state == 2'h1 : _GEN_112; // @[CScratchpad.scala 136:19 138:24]
  wire  _T_13 = auto_mem_out_a_ready & mem_out_a_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_8 = 4'h0 == reqChosen ? 1'h0 : reqIdleBits_0; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_9 = 4'h1 == reqChosen ? 1'h0 : reqIdleBits_1; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_10 = 4'h2 == reqChosen ? 1'h0 : reqIdleBits_2; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_11 = 4'h3 == reqChosen ? 1'h0 : reqIdleBits_3; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_12 = 4'h4 == reqChosen ? 1'h0 : reqIdleBits_4; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_13 = 4'h5 == reqChosen ? 1'h0 : reqIdleBits_5; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_14 = 4'h6 == reqChosen ? 1'h0 : reqIdleBits_6; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_15 = 4'h7 == reqChosen ? 1'h0 : reqIdleBits_7; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_16 = 4'h8 == reqChosen ? 1'h0 : reqIdleBits_8; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_17 = 4'h9 == reqChosen ? 1'h0 : reqIdleBits_9; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_18 = 4'ha == reqChosen ? 1'h0 : reqIdleBits_10; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_19 = 4'hb == reqChosen ? 1'h0 : reqIdleBits_11; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_20 = 4'hc == reqChosen ? 1'h0 : reqIdleBits_12; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_21 = 4'hd == reqChosen ? 1'h0 : reqIdleBits_13; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_22 = 4'he == reqChosen ? 1'h0 : reqIdleBits_14; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_23 = 4'hf == reqChosen ? 1'h0 : reqIdleBits_15; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire [5:0] _GEN_24 = 4'h0 == reqChosen ? totalTx_scratchpadAddress : req_cache_0_scratchpadAddress; // @[CScratchpad.scala 114:30 154:{48,48}]
  wire [5:0] _GEN_25 = 4'h1 == reqChosen ? totalTx_scratchpadAddress : req_cache_1_scratchpadAddress; // @[CScratchpad.scala 114:30 154:{48,48}]
  wire [5:0] _GEN_26 = 4'h2 == reqChosen ? totalTx_scratchpadAddress : req_cache_2_scratchpadAddress; // @[CScratchpad.scala 114:30 154:{48,48}]
  wire [5:0] _GEN_27 = 4'h3 == reqChosen ? totalTx_scratchpadAddress : req_cache_3_scratchpadAddress; // @[CScratchpad.scala 114:30 154:{48,48}]
  wire [5:0] _GEN_28 = 4'h4 == reqChosen ? totalTx_scratchpadAddress : req_cache_4_scratchpadAddress; // @[CScratchpad.scala 114:30 154:{48,48}]
  wire [5:0] _GEN_29 = 4'h5 == reqChosen ? totalTx_scratchpadAddress : req_cache_5_scratchpadAddress; // @[CScratchpad.scala 114:30 154:{48,48}]
  wire [5:0] _GEN_30 = 4'h6 == reqChosen ? totalTx_scratchpadAddress : req_cache_6_scratchpadAddress; // @[CScratchpad.scala 114:30 154:{48,48}]
  wire [5:0] _GEN_31 = 4'h7 == reqChosen ? totalTx_scratchpadAddress : req_cache_7_scratchpadAddress; // @[CScratchpad.scala 114:30 154:{48,48}]
  wire [5:0] _GEN_32 = 4'h8 == reqChosen ? totalTx_scratchpadAddress : req_cache_8_scratchpadAddress; // @[CScratchpad.scala 114:30 154:{48,48}]
  wire [5:0] _GEN_33 = 4'h9 == reqChosen ? totalTx_scratchpadAddress : req_cache_9_scratchpadAddress; // @[CScratchpad.scala 114:30 154:{48,48}]
  wire [5:0] _GEN_34 = 4'ha == reqChosen ? totalTx_scratchpadAddress : req_cache_10_scratchpadAddress; // @[CScratchpad.scala 114:30 154:{48,48}]
  wire [5:0] _GEN_35 = 4'hb == reqChosen ? totalTx_scratchpadAddress : req_cache_11_scratchpadAddress; // @[CScratchpad.scala 114:30 154:{48,48}]
  wire [5:0] _GEN_36 = 4'hc == reqChosen ? totalTx_scratchpadAddress : req_cache_12_scratchpadAddress; // @[CScratchpad.scala 114:30 154:{48,48}]
  wire [5:0] _GEN_37 = 4'hd == reqChosen ? totalTx_scratchpadAddress : req_cache_13_scratchpadAddress; // @[CScratchpad.scala 114:30 154:{48,48}]
  wire [5:0] _GEN_38 = 4'he == reqChosen ? totalTx_scratchpadAddress : req_cache_14_scratchpadAddress; // @[CScratchpad.scala 114:30 154:{48,48}]
  wire [5:0] _GEN_39 = 4'hf == reqChosen ? totalTx_scratchpadAddress : req_cache_15_scratchpadAddress; // @[CScratchpad.scala 114:30 154:{48,48}]
  wire [33:0] _req_cache_memoryLength_T = isBelowLimit ? totalTx_memoryLength : 34'h40; // @[CScratchpad.scala 155:49]
  wire [15:0] _GEN_40 = 4'h0 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_0_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_41 = 4'h1 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_1_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_42 = 4'h2 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_2_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_43 = 4'h3 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_3_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_44 = 4'h4 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_4_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_45 = 4'h5 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_5_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_46 = 4'h6 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_6_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_47 = 4'h7 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_7_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_48 = 4'h8 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_8_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_49 = 4'h9 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_9_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_50 = 4'ha == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_10_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_51 = 4'hb == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_11_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_52 = 4'hc == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_12_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_53 = 4'hd == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_13_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_54 = 4'he == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_14_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_55 = 4'hf == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_15_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [33:0] _totalTx_memoryLength_T_1 = totalTx_memoryLength - 34'h40; // @[CScratchpad.scala 156:54]
  wire [5:0] _totalTx_scratchpadAddress_T_1 = totalTx_scratchpadAddress + 6'h4; // @[CScratchpad.scala 157:64]
  wire [33:0] _totalTx_memoryAddress_T_1 = totalTx_memoryAddress + 34'h40; // @[CScratchpad.scala 158:56]
  wire [1:0] _GEN_56 = isBelowLimit ? 2'h2 : mem_tx_state; // @[CScratchpad.scala 159:28 160:24 102:37]
  wire  _GEN_57 = _T_13 ? _GEN_8 : reqIdleBits_0; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_58 = _T_13 ? _GEN_9 : reqIdleBits_1; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_59 = _T_13 ? _GEN_10 : reqIdleBits_2; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_60 = _T_13 ? _GEN_11 : reqIdleBits_3; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_61 = _T_13 ? _GEN_12 : reqIdleBits_4; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_62 = _T_13 ? _GEN_13 : reqIdleBits_5; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_63 = _T_13 ? _GEN_14 : reqIdleBits_6; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_64 = _T_13 ? _GEN_15 : reqIdleBits_7; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_65 = _T_13 ? _GEN_16 : reqIdleBits_8; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_66 = _T_13 ? _GEN_17 : reqIdleBits_9; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_67 = _T_13 ? _GEN_18 : reqIdleBits_10; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_68 = _T_13 ? _GEN_19 : reqIdleBits_11; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_69 = _T_13 ? _GEN_20 : reqIdleBits_12; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_70 = _T_13 ? _GEN_21 : reqIdleBits_13; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_71 = _T_13 ? _GEN_22 : reqIdleBits_14; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_72 = _T_13 ? _GEN_23 : reqIdleBits_15; // @[CScratchpad.scala 152:28 110:36]
  wire [5:0] _GEN_73 = _T_13 ? _GEN_24 : req_cache_0_scratchpadAddress; // @[CScratchpad.scala 152:28 114:30]
  wire [5:0] _GEN_74 = _T_13 ? _GEN_25 : req_cache_1_scratchpadAddress; // @[CScratchpad.scala 152:28 114:30]
  wire [5:0] _GEN_75 = _T_13 ? _GEN_26 : req_cache_2_scratchpadAddress; // @[CScratchpad.scala 152:28 114:30]
  wire [5:0] _GEN_76 = _T_13 ? _GEN_27 : req_cache_3_scratchpadAddress; // @[CScratchpad.scala 152:28 114:30]
  wire [5:0] _GEN_77 = _T_13 ? _GEN_28 : req_cache_4_scratchpadAddress; // @[CScratchpad.scala 152:28 114:30]
  wire [5:0] _GEN_78 = _T_13 ? _GEN_29 : req_cache_5_scratchpadAddress; // @[CScratchpad.scala 152:28 114:30]
  wire [5:0] _GEN_79 = _T_13 ? _GEN_30 : req_cache_6_scratchpadAddress; // @[CScratchpad.scala 152:28 114:30]
  wire [5:0] _GEN_80 = _T_13 ? _GEN_31 : req_cache_7_scratchpadAddress; // @[CScratchpad.scala 152:28 114:30]
  wire [5:0] _GEN_81 = _T_13 ? _GEN_32 : req_cache_8_scratchpadAddress; // @[CScratchpad.scala 152:28 114:30]
  wire [5:0] _GEN_82 = _T_13 ? _GEN_33 : req_cache_9_scratchpadAddress; // @[CScratchpad.scala 152:28 114:30]
  wire [5:0] _GEN_83 = _T_13 ? _GEN_34 : req_cache_10_scratchpadAddress; // @[CScratchpad.scala 152:28 114:30]
  wire [5:0] _GEN_84 = _T_13 ? _GEN_35 : req_cache_11_scratchpadAddress; // @[CScratchpad.scala 152:28 114:30]
  wire [5:0] _GEN_85 = _T_13 ? _GEN_36 : req_cache_12_scratchpadAddress; // @[CScratchpad.scala 152:28 114:30]
  wire [5:0] _GEN_86 = _T_13 ? _GEN_37 : req_cache_13_scratchpadAddress; // @[CScratchpad.scala 152:28 114:30]
  wire [5:0] _GEN_87 = _T_13 ? _GEN_38 : req_cache_14_scratchpadAddress; // @[CScratchpad.scala 152:28 114:30]
  wire [5:0] _GEN_88 = _T_13 ? _GEN_39 : req_cache_15_scratchpadAddress; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_89 = _T_13 ? _GEN_40 : req_cache_0_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_90 = _T_13 ? _GEN_41 : req_cache_1_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_91 = _T_13 ? _GEN_42 : req_cache_2_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_92 = _T_13 ? _GEN_43 : req_cache_3_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_93 = _T_13 ? _GEN_44 : req_cache_4_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_94 = _T_13 ? _GEN_45 : req_cache_5_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_95 = _T_13 ? _GEN_46 : req_cache_6_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_96 = _T_13 ? _GEN_47 : req_cache_7_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_97 = _T_13 ? _GEN_48 : req_cache_8_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_98 = _T_13 ? _GEN_49 : req_cache_9_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_99 = _T_13 ? _GEN_50 : req_cache_10_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_100 = _T_13 ? _GEN_51 : req_cache_11_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_101 = _T_13 ? _GEN_52 : req_cache_12_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_102 = _T_13 ? _GEN_53 : req_cache_13_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_103 = _T_13 ? _GEN_54 : req_cache_14_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_104 = _T_13 ? _GEN_55 : req_cache_15_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [1:0] _GEN_109 = reqIdleBits_0 & reqIdleBits_1 & reqIdleBits_2 & reqIdleBits_3 & reqIdleBits_4 & reqIdleBits_5 &
    reqIdleBits_6 & reqIdleBits_7 & reqIdleBits_8 & reqIdleBits_9 & reqIdleBits_10 & reqIdleBits_11 & reqIdleBits_12 &
    reqIdleBits_13 & reqIdleBits_14 & reqIdleBits_15 ? 2'h0 : mem_tx_state; // @[CScratchpad.scala 166:40 167:22 102:37]
  wire  _GEN_113 = 2'h1 == mem_tx_state ? _GEN_57 : reqIdleBits_0; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_114 = 2'h1 == mem_tx_state ? _GEN_58 : reqIdleBits_1; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_115 = 2'h1 == mem_tx_state ? _GEN_59 : reqIdleBits_2; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_116 = 2'h1 == mem_tx_state ? _GEN_60 : reqIdleBits_3; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_117 = 2'h1 == mem_tx_state ? _GEN_61 : reqIdleBits_4; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_118 = 2'h1 == mem_tx_state ? _GEN_62 : reqIdleBits_5; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_119 = 2'h1 == mem_tx_state ? _GEN_63 : reqIdleBits_6; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_120 = 2'h1 == mem_tx_state ? _GEN_64 : reqIdleBits_7; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_121 = 2'h1 == mem_tx_state ? _GEN_65 : reqIdleBits_8; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_122 = 2'h1 == mem_tx_state ? _GEN_66 : reqIdleBits_9; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_123 = 2'h1 == mem_tx_state ? _GEN_67 : reqIdleBits_10; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_124 = 2'h1 == mem_tx_state ? _GEN_68 : reqIdleBits_11; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_125 = 2'h1 == mem_tx_state ? _GEN_69 : reqIdleBits_12; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_126 = 2'h1 == mem_tx_state ? _GEN_70 : reqIdleBits_13; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_127 = 2'h1 == mem_tx_state ? _GEN_71 : reqIdleBits_14; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_128 = 2'h1 == mem_tx_state ? _GEN_72 : reqIdleBits_15; // @[CScratchpad.scala 138:24 110:36]
  wire [5:0] _GEN_129 = 2'h1 == mem_tx_state ? _GEN_73 : req_cache_0_scratchpadAddress; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_130 = 2'h1 == mem_tx_state ? _GEN_74 : req_cache_1_scratchpadAddress; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_131 = 2'h1 == mem_tx_state ? _GEN_75 : req_cache_2_scratchpadAddress; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_132 = 2'h1 == mem_tx_state ? _GEN_76 : req_cache_3_scratchpadAddress; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_133 = 2'h1 == mem_tx_state ? _GEN_77 : req_cache_4_scratchpadAddress; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_134 = 2'h1 == mem_tx_state ? _GEN_78 : req_cache_5_scratchpadAddress; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_135 = 2'h1 == mem_tx_state ? _GEN_79 : req_cache_6_scratchpadAddress; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_136 = 2'h1 == mem_tx_state ? _GEN_80 : req_cache_7_scratchpadAddress; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_137 = 2'h1 == mem_tx_state ? _GEN_81 : req_cache_8_scratchpadAddress; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_138 = 2'h1 == mem_tx_state ? _GEN_82 : req_cache_9_scratchpadAddress; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_139 = 2'h1 == mem_tx_state ? _GEN_83 : req_cache_10_scratchpadAddress; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_140 = 2'h1 == mem_tx_state ? _GEN_84 : req_cache_11_scratchpadAddress; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_141 = 2'h1 == mem_tx_state ? _GEN_85 : req_cache_12_scratchpadAddress; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_142 = 2'h1 == mem_tx_state ? _GEN_86 : req_cache_13_scratchpadAddress; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_143 = 2'h1 == mem_tx_state ? _GEN_87 : req_cache_14_scratchpadAddress; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_144 = 2'h1 == mem_tx_state ? _GEN_88 : req_cache_15_scratchpadAddress; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_145 = 2'h1 == mem_tx_state ? _GEN_89 : req_cache_0_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_146 = 2'h1 == mem_tx_state ? _GEN_90 : req_cache_1_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_147 = 2'h1 == mem_tx_state ? _GEN_91 : req_cache_2_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_148 = 2'h1 == mem_tx_state ? _GEN_92 : req_cache_3_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_149 = 2'h1 == mem_tx_state ? _GEN_93 : req_cache_4_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_150 = 2'h1 == mem_tx_state ? _GEN_94 : req_cache_5_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_151 = 2'h1 == mem_tx_state ? _GEN_95 : req_cache_6_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_152 = 2'h1 == mem_tx_state ? _GEN_96 : req_cache_7_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_153 = 2'h1 == mem_tx_state ? _GEN_97 : req_cache_8_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_154 = 2'h1 == mem_tx_state ? _GEN_98 : req_cache_9_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_155 = 2'h1 == mem_tx_state ? _GEN_99 : req_cache_10_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_156 = 2'h1 == mem_tx_state ? _GEN_100 : req_cache_11_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_157 = 2'h1 == mem_tx_state ? _GEN_101 : req_cache_12_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_158 = 2'h1 == mem_tx_state ? _GEN_102 : req_cache_13_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_159 = 2'h1 == mem_tx_state ? _GEN_103 : req_cache_14_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_160 = 2'h1 == mem_tx_state ? _GEN_104 : req_cache_15_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire  _GEN_171 = 2'h0 == mem_tx_state ? reqIdleBits_0 : _GEN_113; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_172 = 2'h0 == mem_tx_state ? reqIdleBits_1 : _GEN_114; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_173 = 2'h0 == mem_tx_state ? reqIdleBits_2 : _GEN_115; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_174 = 2'h0 == mem_tx_state ? reqIdleBits_3 : _GEN_116; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_175 = 2'h0 == mem_tx_state ? reqIdleBits_4 : _GEN_117; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_176 = 2'h0 == mem_tx_state ? reqIdleBits_5 : _GEN_118; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_177 = 2'h0 == mem_tx_state ? reqIdleBits_6 : _GEN_119; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_178 = 2'h0 == mem_tx_state ? reqIdleBits_7 : _GEN_120; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_179 = 2'h0 == mem_tx_state ? reqIdleBits_8 : _GEN_121; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_180 = 2'h0 == mem_tx_state ? reqIdleBits_9 : _GEN_122; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_181 = 2'h0 == mem_tx_state ? reqIdleBits_10 : _GEN_123; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_182 = 2'h0 == mem_tx_state ? reqIdleBits_11 : _GEN_124; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_183 = 2'h0 == mem_tx_state ? reqIdleBits_12 : _GEN_125; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_184 = 2'h0 == mem_tx_state ? reqIdleBits_13 : _GEN_126; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_185 = 2'h0 == mem_tx_state ? reqIdleBits_14 : _GEN_127; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_186 = 2'h0 == mem_tx_state ? reqIdleBits_15 : _GEN_128; // @[CScratchpad.scala 138:24 110:36]
  wire [5:0] _GEN_187 = 2'h0 == mem_tx_state ? req_cache_0_scratchpadAddress : _GEN_129; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_188 = 2'h0 == mem_tx_state ? req_cache_1_scratchpadAddress : _GEN_130; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_189 = 2'h0 == mem_tx_state ? req_cache_2_scratchpadAddress : _GEN_131; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_190 = 2'h0 == mem_tx_state ? req_cache_3_scratchpadAddress : _GEN_132; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_191 = 2'h0 == mem_tx_state ? req_cache_4_scratchpadAddress : _GEN_133; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_192 = 2'h0 == mem_tx_state ? req_cache_5_scratchpadAddress : _GEN_134; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_193 = 2'h0 == mem_tx_state ? req_cache_6_scratchpadAddress : _GEN_135; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_194 = 2'h0 == mem_tx_state ? req_cache_7_scratchpadAddress : _GEN_136; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_195 = 2'h0 == mem_tx_state ? req_cache_8_scratchpadAddress : _GEN_137; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_196 = 2'h0 == mem_tx_state ? req_cache_9_scratchpadAddress : _GEN_138; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_197 = 2'h0 == mem_tx_state ? req_cache_10_scratchpadAddress : _GEN_139; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_198 = 2'h0 == mem_tx_state ? req_cache_11_scratchpadAddress : _GEN_140; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_199 = 2'h0 == mem_tx_state ? req_cache_12_scratchpadAddress : _GEN_141; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_200 = 2'h0 == mem_tx_state ? req_cache_13_scratchpadAddress : _GEN_142; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_201 = 2'h0 == mem_tx_state ? req_cache_14_scratchpadAddress : _GEN_143; // @[CScratchpad.scala 138:24 114:30]
  wire [5:0] _GEN_202 = 2'h0 == mem_tx_state ? req_cache_15_scratchpadAddress : _GEN_144; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_203 = 2'h0 == mem_tx_state ? req_cache_0_memoryLength : _GEN_145; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_204 = 2'h0 == mem_tx_state ? req_cache_1_memoryLength : _GEN_146; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_205 = 2'h0 == mem_tx_state ? req_cache_2_memoryLength : _GEN_147; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_206 = 2'h0 == mem_tx_state ? req_cache_3_memoryLength : _GEN_148; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_207 = 2'h0 == mem_tx_state ? req_cache_4_memoryLength : _GEN_149; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_208 = 2'h0 == mem_tx_state ? req_cache_5_memoryLength : _GEN_150; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_209 = 2'h0 == mem_tx_state ? req_cache_6_memoryLength : _GEN_151; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_210 = 2'h0 == mem_tx_state ? req_cache_7_memoryLength : _GEN_152; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_211 = 2'h0 == mem_tx_state ? req_cache_8_memoryLength : _GEN_153; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_212 = 2'h0 == mem_tx_state ? req_cache_9_memoryLength : _GEN_154; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_213 = 2'h0 == mem_tx_state ? req_cache_10_memoryLength : _GEN_155; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_214 = 2'h0 == mem_tx_state ? req_cache_11_memoryLength : _GEN_156; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_215 = 2'h0 == mem_tx_state ? req_cache_12_memoryLength : _GEN_157; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_216 = 2'h0 == mem_tx_state ? req_cache_13_memoryLength : _GEN_158; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_217 = 2'h0 == mem_tx_state ? req_cache_14_memoryLength : _GEN_159; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_218 = 2'h0 == mem_tx_state ? req_cache_15_memoryLength : _GEN_160; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_220 = 4'h1 == auto_mem_out_d_bits_source ? req_cache_1_memoryLength : req_cache_0_memoryLength; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_221 = 4'h2 == auto_mem_out_d_bits_source ? req_cache_2_memoryLength : _GEN_220; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_222 = 4'h3 == auto_mem_out_d_bits_source ? req_cache_3_memoryLength : _GEN_221; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_223 = 4'h4 == auto_mem_out_d_bits_source ? req_cache_4_memoryLength : _GEN_222; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_224 = 4'h5 == auto_mem_out_d_bits_source ? req_cache_5_memoryLength : _GEN_223; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_225 = 4'h6 == auto_mem_out_d_bits_source ? req_cache_6_memoryLength : _GEN_224; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_226 = 4'h7 == auto_mem_out_d_bits_source ? req_cache_7_memoryLength : _GEN_225; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_227 = 4'h8 == auto_mem_out_d_bits_source ? req_cache_8_memoryLength : _GEN_226; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_228 = 4'h9 == auto_mem_out_d_bits_source ? req_cache_9_memoryLength : _GEN_227; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_229 = 4'ha == auto_mem_out_d_bits_source ? req_cache_10_memoryLength : _GEN_228; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_230 = 4'hb == auto_mem_out_d_bits_source ? req_cache_11_memoryLength : _GEN_229; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_231 = 4'hc == auto_mem_out_d_bits_source ? req_cache_12_memoryLength : _GEN_230; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_232 = 4'hd == auto_mem_out_d_bits_source ? req_cache_13_memoryLength : _GEN_231; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_233 = 4'he == auto_mem_out_d_bits_source ? req_cache_14_memoryLength : _GEN_232; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_234 = 4'hf == auto_mem_out_d_bits_source ? req_cache_15_memoryLength : _GEN_233; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_235 = _GEN_234 >= 16'h40 ? 16'h40 : _GEN_234; // @[CScratchpad.scala 174:55 175:39 177:39]
  wire [5:0] _GEN_237 = 4'h1 == auto_mem_out_d_bits_source ? req_cache_1_scratchpadAddress :
    req_cache_0_scratchpadAddress; // @[CScratchpad.scala 179:{41,41}]
  wire [5:0] _GEN_238 = 4'h2 == auto_mem_out_d_bits_source ? req_cache_2_scratchpadAddress : _GEN_237; // @[CScratchpad.scala 179:{41,41}]
  wire [5:0] _GEN_239 = 4'h3 == auto_mem_out_d_bits_source ? req_cache_3_scratchpadAddress : _GEN_238; // @[CScratchpad.scala 179:{41,41}]
  wire [5:0] _GEN_240 = 4'h4 == auto_mem_out_d_bits_source ? req_cache_4_scratchpadAddress : _GEN_239; // @[CScratchpad.scala 179:{41,41}]
  wire [5:0] _GEN_241 = 4'h5 == auto_mem_out_d_bits_source ? req_cache_5_scratchpadAddress : _GEN_240; // @[CScratchpad.scala 179:{41,41}]
  wire [5:0] _GEN_242 = 4'h6 == auto_mem_out_d_bits_source ? req_cache_6_scratchpadAddress : _GEN_241; // @[CScratchpad.scala 179:{41,41}]
  wire [5:0] _GEN_243 = 4'h7 == auto_mem_out_d_bits_source ? req_cache_7_scratchpadAddress : _GEN_242; // @[CScratchpad.scala 179:{41,41}]
  wire [5:0] _GEN_244 = 4'h8 == auto_mem_out_d_bits_source ? req_cache_8_scratchpadAddress : _GEN_243; // @[CScratchpad.scala 179:{41,41}]
  wire [5:0] _GEN_245 = 4'h9 == auto_mem_out_d_bits_source ? req_cache_9_scratchpadAddress : _GEN_244; // @[CScratchpad.scala 179:{41,41}]
  wire [5:0] _GEN_246 = 4'ha == auto_mem_out_d_bits_source ? req_cache_10_scratchpadAddress : _GEN_245; // @[CScratchpad.scala 179:{41,41}]
  wire [5:0] _GEN_247 = 4'hb == auto_mem_out_d_bits_source ? req_cache_11_scratchpadAddress : _GEN_246; // @[CScratchpad.scala 179:{41,41}]
  wire [5:0] _GEN_248 = 4'hc == auto_mem_out_d_bits_source ? req_cache_12_scratchpadAddress : _GEN_247; // @[CScratchpad.scala 179:{41,41}]
  wire [5:0] _GEN_249 = 4'hd == auto_mem_out_d_bits_source ? req_cache_13_scratchpadAddress : _GEN_248; // @[CScratchpad.scala 179:{41,41}]
  wire [5:0] _GEN_250 = 4'he == auto_mem_out_d_bits_source ? req_cache_14_scratchpadAddress : _GEN_249; // @[CScratchpad.scala 179:{41,41}]
  wire [5:0] _GEN_251 = 4'hf == auto_mem_out_d_bits_source ? req_cache_15_scratchpadAddress : _GEN_250; // @[CScratchpad.scala 179:{41,41}]
  wire  _T_31 = loader_io_cache_block_in_ready & loader_io_cache_block_in_valid; // @[Decoupled.scala 51:35]
  wire [5:0] _req_cache_scratchpadAddress_T_1 = _GEN_251 + 6'h4; // @[CScratchpad.scala 183:82]
  wire  mem_out_d_ready = loader_io_cache_block_in_ready; // @[Nodes.scala 1212:84 CScratchpad.scala 180:19]
  wire  _T_36 = mem_out_d_ready & auto_mem_out_d_valid; // @[Decoupled.scala 51:35]
  wire [15:0] _req_cache_memoryLength_T_2 = _GEN_234 - 16'h40; // @[CScratchpad.scala 210:72]
  wire  _GEN_445 = 4'h0 == auto_mem_out_d_bits_source | _GEN_171; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_446 = 4'h1 == auto_mem_out_d_bits_source | _GEN_172; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_447 = 4'h2 == auto_mem_out_d_bits_source | _GEN_173; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_448 = 4'h3 == auto_mem_out_d_bits_source | _GEN_174; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_449 = 4'h4 == auto_mem_out_d_bits_source | _GEN_175; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_450 = 4'h5 == auto_mem_out_d_bits_source | _GEN_176; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_451 = 4'h6 == auto_mem_out_d_bits_source | _GEN_177; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_452 = 4'h7 == auto_mem_out_d_bits_source | _GEN_178; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_453 = 4'h8 == auto_mem_out_d_bits_source | _GEN_179; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_454 = 4'h9 == auto_mem_out_d_bits_source | _GEN_180; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_455 = 4'ha == auto_mem_out_d_bits_source | _GEN_181; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_456 = 4'hb == auto_mem_out_d_bits_source | _GEN_182; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_457 = 4'hc == auto_mem_out_d_bits_source | _GEN_183; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_458 = 4'hd == auto_mem_out_d_bits_source | _GEN_184; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_459 = 4'he == auto_mem_out_d_bits_source | _GEN_185; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_460 = 4'hf == auto_mem_out_d_bits_source | _GEN_186; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_461 = _GEN_234 <= 16'h40 ? _GEN_445 : _GEN_171; // @[CScratchpad.scala 212:57]
  wire  _GEN_462 = _GEN_234 <= 16'h40 ? _GEN_446 : _GEN_172; // @[CScratchpad.scala 212:57]
  wire  _GEN_463 = _GEN_234 <= 16'h40 ? _GEN_447 : _GEN_173; // @[CScratchpad.scala 212:57]
  wire  _GEN_464 = _GEN_234 <= 16'h40 ? _GEN_448 : _GEN_174; // @[CScratchpad.scala 212:57]
  wire  _GEN_465 = _GEN_234 <= 16'h40 ? _GEN_449 : _GEN_175; // @[CScratchpad.scala 212:57]
  wire  _GEN_466 = _GEN_234 <= 16'h40 ? _GEN_450 : _GEN_176; // @[CScratchpad.scala 212:57]
  wire  _GEN_467 = _GEN_234 <= 16'h40 ? _GEN_451 : _GEN_177; // @[CScratchpad.scala 212:57]
  wire  _GEN_468 = _GEN_234 <= 16'h40 ? _GEN_452 : _GEN_178; // @[CScratchpad.scala 212:57]
  wire  _GEN_469 = _GEN_234 <= 16'h40 ? _GEN_453 : _GEN_179; // @[CScratchpad.scala 212:57]
  wire  _GEN_470 = _GEN_234 <= 16'h40 ? _GEN_454 : _GEN_180; // @[CScratchpad.scala 212:57]
  wire  _GEN_471 = _GEN_234 <= 16'h40 ? _GEN_455 : _GEN_181; // @[CScratchpad.scala 212:57]
  wire  _GEN_472 = _GEN_234 <= 16'h40 ? _GEN_456 : _GEN_182; // @[CScratchpad.scala 212:57]
  wire  _GEN_473 = _GEN_234 <= 16'h40 ? _GEN_457 : _GEN_183; // @[CScratchpad.scala 212:57]
  wire  _GEN_474 = _GEN_234 <= 16'h40 ? _GEN_458 : _GEN_184; // @[CScratchpad.scala 212:57]
  wire  _GEN_475 = _GEN_234 <= 16'h40 ? _GEN_459 : _GEN_185; // @[CScratchpad.scala 212:57]
  wire  _GEN_476 = _GEN_234 <= 16'h40 ? _GEN_460 : _GEN_186; // @[CScratchpad.scala 212:57]
  wire  _GEN_494 = _T_36 ? _GEN_461 : _GEN_171; // @[CScratchpad.scala 209:24]
  wire  _GEN_495 = _T_36 ? _GEN_462 : _GEN_172; // @[CScratchpad.scala 209:24]
  wire  _GEN_496 = _T_36 ? _GEN_463 : _GEN_173; // @[CScratchpad.scala 209:24]
  wire  _GEN_497 = _T_36 ? _GEN_464 : _GEN_174; // @[CScratchpad.scala 209:24]
  wire  _GEN_498 = _T_36 ? _GEN_465 : _GEN_175; // @[CScratchpad.scala 209:24]
  wire  _GEN_499 = _T_36 ? _GEN_466 : _GEN_176; // @[CScratchpad.scala 209:24]
  wire  _GEN_500 = _T_36 ? _GEN_467 : _GEN_177; // @[CScratchpad.scala 209:24]
  wire  _GEN_501 = _T_36 ? _GEN_468 : _GEN_178; // @[CScratchpad.scala 209:24]
  wire  _GEN_502 = _T_36 ? _GEN_469 : _GEN_179; // @[CScratchpad.scala 209:24]
  wire  _GEN_503 = _T_36 ? _GEN_470 : _GEN_180; // @[CScratchpad.scala 209:24]
  wire  _GEN_504 = _T_36 ? _GEN_471 : _GEN_181; // @[CScratchpad.scala 209:24]
  wire  _GEN_505 = _T_36 ? _GEN_472 : _GEN_182; // @[CScratchpad.scala 209:24]
  wire  _GEN_506 = _T_36 ? _GEN_473 : _GEN_183; // @[CScratchpad.scala 209:24]
  wire  _GEN_507 = _T_36 ? _GEN_474 : _GEN_184; // @[CScratchpad.scala 209:24]
  wire  _GEN_508 = _T_36 ? _GEN_475 : _GEN_185; // @[CScratchpad.scala 209:24]
  wire  _GEN_509 = _T_36 ? _GEN_476 : _GEN_186; // @[CScratchpad.scala 209:24]
  CScratchpadPackedSubwordLoader loader ( // @[CScratchpad.scala 94:30]
    .clock(loader_clock),
    .reset(loader_reset),
    .io_cache_block_in_ready(loader_io_cache_block_in_ready),
    .io_cache_block_in_valid(loader_io_cache_block_in_valid),
    .io_cache_block_in_bits_dat(loader_io_cache_block_in_bits_dat),
    .io_cache_block_in_bits_len(loader_io_cache_block_in_bits_len),
    .io_cache_block_in_bits_idxBase(loader_io_cache_block_in_bits_idxBase),
    .io_sp_write_out_valid(loader_io_sp_write_out_valid),
    .io_sp_write_out_bits_dat(loader_io_sp_write_out_bits_dat),
    .io_sp_write_out_bits_idx(loader_io_sp_write_out_bits_idx)
  );
  assign mem_rval_en = mem_rval_en_pipe_0;
  assign mem_rval_addr = mem_rval_addr_pipe_0;
  assign mem_rval_data = mem[mem_rval_addr]; // @[CScratchpad.scala 92:24]
  assign mem_MPORT_data = loader_io_sp_write_out_bits_dat;
  assign mem_MPORT_addr = loader_io_sp_write_out_bits_idx;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = loader_io_sp_write_out_valid;
  assign mem_MPORT_1_data = 128'h0;
  assign mem_MPORT_1_addr = 6'h0;
  assign mem_MPORT_1_mask = 1'h1;
  assign mem_MPORT_1_en = 1'h0;
  assign auto_mem_out_a_valid = 2'h0 == mem_tx_state ? mem_tx_state == 2'h1 : _GEN_112; // @[CScratchpad.scala 136:19 138:24]
  assign auto_mem_out_a_bits_size = txEmitLengthLg[2:0]; // @[Edges.scala 447:17 450:15]
  assign auto_mem_out_a_bits_source = reqIdleBits_0 ? 4'h0 : _reqChosen_T_13; // @[Mux.scala 47:70]
  assign auto_mem_out_a_bits_address = totalTx_memoryAddress; // @[Edges.scala 447:17 452:15]
  assign auto_mem_out_a_bits_mask = {x1_a_bits_a_mask_hi,x1_a_bits_a_mask_lo}; // @[Cat.scala 33:92]
  assign auto_mem_out_d_ready = loader_io_cache_block_in_ready; // @[Nodes.scala 1212:84 CScratchpad.scala 180:19]
  assign access_readRes_valid = access_readRes_valid_REG; // @[CScratchpad.scala 103:24]
  assign access_readRes_bits = mem_rval_data; // @[CScratchpad.scala 105:23]
  assign loader_clock = clock;
  assign loader_reset = reset;
  assign loader_io_cache_block_in_valid = auto_mem_out_d_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign loader_io_cache_block_in_bits_dat = auto_mem_out_d_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign loader_io_cache_block_in_bits_len = _GEN_235[6:0];
  assign loader_io_cache_block_in_bits_idxBase = 4'hf == auto_mem_out_d_bits_source ? req_cache_15_scratchpadAddress :
    _GEN_250; // @[CScratchpad.scala 179:{41,41}]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[CScratchpad.scala 92:24]
    end
    if (mem_MPORT_1_en & mem_MPORT_1_mask) begin
      mem[mem_MPORT_1_addr] <= mem_MPORT_1_data; // @[CScratchpad.scala 92:24]
    end
    mem_rval_en_pipe_0 <= access_readReq_valid;
    if (access_readReq_valid) begin
      mem_rval_addr_pipe_0 <= 6'h0;
    end
    if (reset) begin // @[CScratchpad.scala 102:37]
      mem_tx_state <= 2'h0; // @[CScratchpad.scala 102:37]
    end else if (!(2'h0 == mem_tx_state)) begin // @[CScratchpad.scala 138:24]
      if (2'h1 == mem_tx_state) begin // @[CScratchpad.scala 138:24]
        if (_T_13) begin // @[CScratchpad.scala 152:28]
          mem_tx_state <= _GEN_56;
        end
      end else if (2'h2 == mem_tx_state) begin // @[CScratchpad.scala 138:24]
        mem_tx_state <= _GEN_109;
      end
    end
    access_readRes_valid_REG <= access_readReq_valid; // @[CScratchpad.scala 85:30]
    reqIdleBits_0 <= reset | _GEN_494; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_1 <= reset | _GEN_495; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_2 <= reset | _GEN_496; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_3 <= reset | _GEN_497; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_4 <= reset | _GEN_498; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_5 <= reset | _GEN_499; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_6 <= reset | _GEN_500; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_7 <= reset | _GEN_501; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_8 <= reset | _GEN_502; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_9 <= reset | _GEN_503; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_10 <= reset | _GEN_504; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_11 <= reset | _GEN_505; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_12 <= reset | _GEN_506; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_13 <= reset | _GEN_507; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_14 <= reset | _GEN_508; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_15 <= reset | _GEN_509; // @[CScratchpad.scala 110:{36,36}]
    if (_T_31) begin // @[CScratchpad.scala 182:39]
      if (4'h0 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 183:42]
        req_cache_0_scratchpadAddress <= _req_cache_scratchpadAddress_T_1; // @[CScratchpad.scala 183:42]
      end else begin
        req_cache_0_scratchpadAddress <= _GEN_187;
      end
    end else begin
      req_cache_0_scratchpadAddress <= _GEN_187;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h0 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_0_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_0_memoryLength <= _GEN_203;
      end
    end else begin
      req_cache_0_memoryLength <= _GEN_203;
    end
    if (_T_31) begin // @[CScratchpad.scala 182:39]
      if (4'h1 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 183:42]
        req_cache_1_scratchpadAddress <= _req_cache_scratchpadAddress_T_1; // @[CScratchpad.scala 183:42]
      end else begin
        req_cache_1_scratchpadAddress <= _GEN_188;
      end
    end else begin
      req_cache_1_scratchpadAddress <= _GEN_188;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h1 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_1_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_1_memoryLength <= _GEN_204;
      end
    end else begin
      req_cache_1_memoryLength <= _GEN_204;
    end
    if (_T_31) begin // @[CScratchpad.scala 182:39]
      if (4'h2 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 183:42]
        req_cache_2_scratchpadAddress <= _req_cache_scratchpadAddress_T_1; // @[CScratchpad.scala 183:42]
      end else begin
        req_cache_2_scratchpadAddress <= _GEN_189;
      end
    end else begin
      req_cache_2_scratchpadAddress <= _GEN_189;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h2 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_2_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_2_memoryLength <= _GEN_205;
      end
    end else begin
      req_cache_2_memoryLength <= _GEN_205;
    end
    if (_T_31) begin // @[CScratchpad.scala 182:39]
      if (4'h3 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 183:42]
        req_cache_3_scratchpadAddress <= _req_cache_scratchpadAddress_T_1; // @[CScratchpad.scala 183:42]
      end else begin
        req_cache_3_scratchpadAddress <= _GEN_190;
      end
    end else begin
      req_cache_3_scratchpadAddress <= _GEN_190;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h3 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_3_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_3_memoryLength <= _GEN_206;
      end
    end else begin
      req_cache_3_memoryLength <= _GEN_206;
    end
    if (_T_31) begin // @[CScratchpad.scala 182:39]
      if (4'h4 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 183:42]
        req_cache_4_scratchpadAddress <= _req_cache_scratchpadAddress_T_1; // @[CScratchpad.scala 183:42]
      end else begin
        req_cache_4_scratchpadAddress <= _GEN_191;
      end
    end else begin
      req_cache_4_scratchpadAddress <= _GEN_191;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h4 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_4_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_4_memoryLength <= _GEN_207;
      end
    end else begin
      req_cache_4_memoryLength <= _GEN_207;
    end
    if (_T_31) begin // @[CScratchpad.scala 182:39]
      if (4'h5 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 183:42]
        req_cache_5_scratchpadAddress <= _req_cache_scratchpadAddress_T_1; // @[CScratchpad.scala 183:42]
      end else begin
        req_cache_5_scratchpadAddress <= _GEN_192;
      end
    end else begin
      req_cache_5_scratchpadAddress <= _GEN_192;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h5 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_5_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_5_memoryLength <= _GEN_208;
      end
    end else begin
      req_cache_5_memoryLength <= _GEN_208;
    end
    if (_T_31) begin // @[CScratchpad.scala 182:39]
      if (4'h6 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 183:42]
        req_cache_6_scratchpadAddress <= _req_cache_scratchpadAddress_T_1; // @[CScratchpad.scala 183:42]
      end else begin
        req_cache_6_scratchpadAddress <= _GEN_193;
      end
    end else begin
      req_cache_6_scratchpadAddress <= _GEN_193;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h6 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_6_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_6_memoryLength <= _GEN_209;
      end
    end else begin
      req_cache_6_memoryLength <= _GEN_209;
    end
    if (_T_31) begin // @[CScratchpad.scala 182:39]
      if (4'h7 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 183:42]
        req_cache_7_scratchpadAddress <= _req_cache_scratchpadAddress_T_1; // @[CScratchpad.scala 183:42]
      end else begin
        req_cache_7_scratchpadAddress <= _GEN_194;
      end
    end else begin
      req_cache_7_scratchpadAddress <= _GEN_194;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h7 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_7_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_7_memoryLength <= _GEN_210;
      end
    end else begin
      req_cache_7_memoryLength <= _GEN_210;
    end
    if (_T_31) begin // @[CScratchpad.scala 182:39]
      if (4'h8 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 183:42]
        req_cache_8_scratchpadAddress <= _req_cache_scratchpadAddress_T_1; // @[CScratchpad.scala 183:42]
      end else begin
        req_cache_8_scratchpadAddress <= _GEN_195;
      end
    end else begin
      req_cache_8_scratchpadAddress <= _GEN_195;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h8 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_8_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_8_memoryLength <= _GEN_211;
      end
    end else begin
      req_cache_8_memoryLength <= _GEN_211;
    end
    if (_T_31) begin // @[CScratchpad.scala 182:39]
      if (4'h9 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 183:42]
        req_cache_9_scratchpadAddress <= _req_cache_scratchpadAddress_T_1; // @[CScratchpad.scala 183:42]
      end else begin
        req_cache_9_scratchpadAddress <= _GEN_196;
      end
    end else begin
      req_cache_9_scratchpadAddress <= _GEN_196;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h9 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_9_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_9_memoryLength <= _GEN_212;
      end
    end else begin
      req_cache_9_memoryLength <= _GEN_212;
    end
    if (_T_31) begin // @[CScratchpad.scala 182:39]
      if (4'ha == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 183:42]
        req_cache_10_scratchpadAddress <= _req_cache_scratchpadAddress_T_1; // @[CScratchpad.scala 183:42]
      end else begin
        req_cache_10_scratchpadAddress <= _GEN_197;
      end
    end else begin
      req_cache_10_scratchpadAddress <= _GEN_197;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'ha == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_10_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_10_memoryLength <= _GEN_213;
      end
    end else begin
      req_cache_10_memoryLength <= _GEN_213;
    end
    if (_T_31) begin // @[CScratchpad.scala 182:39]
      if (4'hb == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 183:42]
        req_cache_11_scratchpadAddress <= _req_cache_scratchpadAddress_T_1; // @[CScratchpad.scala 183:42]
      end else begin
        req_cache_11_scratchpadAddress <= _GEN_198;
      end
    end else begin
      req_cache_11_scratchpadAddress <= _GEN_198;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'hb == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_11_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_11_memoryLength <= _GEN_214;
      end
    end else begin
      req_cache_11_memoryLength <= _GEN_214;
    end
    if (_T_31) begin // @[CScratchpad.scala 182:39]
      if (4'hc == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 183:42]
        req_cache_12_scratchpadAddress <= _req_cache_scratchpadAddress_T_1; // @[CScratchpad.scala 183:42]
      end else begin
        req_cache_12_scratchpadAddress <= _GEN_199;
      end
    end else begin
      req_cache_12_scratchpadAddress <= _GEN_199;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'hc == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_12_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_12_memoryLength <= _GEN_215;
      end
    end else begin
      req_cache_12_memoryLength <= _GEN_215;
    end
    if (_T_31) begin // @[CScratchpad.scala 182:39]
      if (4'hd == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 183:42]
        req_cache_13_scratchpadAddress <= _req_cache_scratchpadAddress_T_1; // @[CScratchpad.scala 183:42]
      end else begin
        req_cache_13_scratchpadAddress <= _GEN_200;
      end
    end else begin
      req_cache_13_scratchpadAddress <= _GEN_200;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'hd == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_13_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_13_memoryLength <= _GEN_216;
      end
    end else begin
      req_cache_13_memoryLength <= _GEN_216;
    end
    if (_T_31) begin // @[CScratchpad.scala 182:39]
      if (4'he == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 183:42]
        req_cache_14_scratchpadAddress <= _req_cache_scratchpadAddress_T_1; // @[CScratchpad.scala 183:42]
      end else begin
        req_cache_14_scratchpadAddress <= _GEN_201;
      end
    end else begin
      req_cache_14_scratchpadAddress <= _GEN_201;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'he == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_14_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_14_memoryLength <= _GEN_217;
      end
    end else begin
      req_cache_14_memoryLength <= _GEN_217;
    end
    if (_T_31) begin // @[CScratchpad.scala 182:39]
      if (4'hf == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 183:42]
        req_cache_15_scratchpadAddress <= _req_cache_scratchpadAddress_T_1; // @[CScratchpad.scala 183:42]
      end else begin
        req_cache_15_scratchpadAddress <= _GEN_202;
      end
    end else begin
      req_cache_15_scratchpadAddress <= _GEN_202;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'hf == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_15_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_15_memoryLength <= _GEN_218;
      end
    end else begin
      req_cache_15_memoryLength <= _GEN_218;
    end
    if (!(2'h0 == mem_tx_state)) begin // @[CScratchpad.scala 138:24]
      if (2'h1 == mem_tx_state) begin // @[CScratchpad.scala 138:24]
        if (_T_13) begin // @[CScratchpad.scala 152:28]
          totalTx_memoryAddress <= _totalTx_memoryAddress_T_1; // @[CScratchpad.scala 158:31]
        end
      end
    end
    if (!(2'h0 == mem_tx_state)) begin // @[CScratchpad.scala 138:24]
      if (2'h1 == mem_tx_state) begin // @[CScratchpad.scala 138:24]
        if (_T_13) begin // @[CScratchpad.scala 152:28]
          totalTx_scratchpadAddress <= _totalTx_scratchpadAddress_T_1; // @[CScratchpad.scala 157:35]
        end
      end
    end
    if (!(2'h0 == mem_tx_state)) begin // @[CScratchpad.scala 138:24]
      if (2'h1 == mem_tx_state) begin // @[CScratchpad.scala 138:24]
        if (_T_13) begin // @[CScratchpad.scala 152:28]
          totalTx_memoryLength <= _totalTx_memoryLength_T_1; // @[CScratchpad.scala 156:30]
        end
      end
    end
  end
endmodule
module CScratchpadPackedSubwordLoader_1(
  input        clock,
  input        reset,
  output       io_cache_block_in_ready,
  input        io_cache_block_in_valid,
  input  [6:0] io_cache_block_in_bits_len,
  output       io_sp_write_out_valid
);
  reg [6:0] lenRemainingFromReq; // @[CScratchpadPackedSubwordLoader.scala 18:32]
  reg  state; // @[CScratchpadPackedSubwordLoader.scala 21:22]
  wire  _io_cache_block_in_ready_T = ~state; // @[CScratchpadPackedSubwordLoader.scala 22:36]
  wire  _T_1 = io_cache_block_in_ready & io_cache_block_in_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_0 = _T_1 | state; // @[CScratchpadPackedSubwordLoader.scala 34:36 35:15 21:22]
  wire [6:0] _lenRemainingFromReq_T_1 = lenRemainingFromReq - 7'h20; // @[CScratchpadPackedSubwordLoader.scala 53:54]
  wire  _GEN_6 = lenRemainingFromReq == 7'h20 ? 1'h0 : state; // @[CScratchpadPackedSubwordLoader.scala 54:60 55:19 21:22]
  assign io_cache_block_in_ready = ~state; // @[CScratchpadPackedSubwordLoader.scala 22:36]
  assign io_sp_write_out_valid = _io_cache_block_in_ready_T ? 1'h0 : state; // @[CScratchpadPackedSubwordLoader.scala 32:17 24:25]
  always @(posedge clock) begin
    if (_io_cache_block_in_ready_T) begin // @[CScratchpadPackedSubwordLoader.scala 32:17]
      if (_T_1) begin // @[CScratchpadPackedSubwordLoader.scala 34:36]
        lenRemainingFromReq <= io_cache_block_in_bits_len; // @[CScratchpadPackedSubwordLoader.scala 38:29]
      end
    end else if (state) begin // @[CScratchpadPackedSubwordLoader.scala 32:17]
      if (io_sp_write_out_valid) begin // @[CScratchpadPackedSubwordLoader.scala 48:34]
        lenRemainingFromReq <= _lenRemainingFromReq_T_1;
      end
    end
    if (reset) begin // @[CScratchpadPackedSubwordLoader.scala 21:22]
      state <= 1'h0; // @[CScratchpadPackedSubwordLoader.scala 21:22]
    end else if (_io_cache_block_in_ready_T) begin // @[CScratchpadPackedSubwordLoader.scala 32:17]
      state <= _GEN_0;
    end else if (state) begin // @[CScratchpadPackedSubwordLoader.scala 32:17]
      if (io_sp_write_out_valid) begin // @[CScratchpadPackedSubwordLoader.scala 48:34]
        state <= _GEN_6;
      end
    end
  end
endmodule
module CScratchpad_1(
  input         clock,
  input         reset,
  input         auto_mem_out_a_ready,
  output        auto_mem_out_a_valid,
  output [2:0]  auto_mem_out_a_bits_size,
  output [3:0]  auto_mem_out_a_bits_source,
  output [33:0] auto_mem_out_a_bits_address,
  output [63:0] auto_mem_out_a_bits_mask,
  output        auto_mem_out_d_ready,
  input         auto_mem_out_d_valid,
  input  [3:0]  auto_mem_out_d_bits_source
);
  wire  loader_clock; // @[CScratchpad.scala 94:30]
  wire  loader_reset; // @[CScratchpad.scala 94:30]
  wire  loader_io_cache_block_in_ready; // @[CScratchpad.scala 94:30]
  wire  loader_io_cache_block_in_valid; // @[CScratchpad.scala 94:30]
  wire [6:0] loader_io_cache_block_in_bits_len; // @[CScratchpad.scala 94:30]
  wire  loader_io_sp_write_out_valid; // @[CScratchpad.scala 94:30]
  reg [1:0] mem_tx_state; // @[CScratchpad.scala 102:37]
  reg  reqIdleBits_0; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_1; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_2; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_3; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_4; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_5; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_6; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_7; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_8; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_9; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_10; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_11; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_12; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_13; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_14; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_15; // @[CScratchpad.scala 110:36]
  wire  reqAvailable = reqIdleBits_0 | reqIdleBits_1 | reqIdleBits_2 | reqIdleBits_3 | reqIdleBits_4 | reqIdleBits_5 |
    reqIdleBits_6 | reqIdleBits_7 | reqIdleBits_8 | reqIdleBits_9 | reqIdleBits_10 | reqIdleBits_11 | reqIdleBits_12 |
    reqIdleBits_13 | reqIdleBits_14 | reqIdleBits_15; // @[CScratchpad.scala 111:51]
  wire [3:0] _reqChosen_T = reqIdleBits_14 ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_1 = reqIdleBits_13 ? 4'hd : _reqChosen_T; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_2 = reqIdleBits_12 ? 4'hc : _reqChosen_T_1; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_3 = reqIdleBits_11 ? 4'hb : _reqChosen_T_2; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_4 = reqIdleBits_10 ? 4'ha : _reqChosen_T_3; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_5 = reqIdleBits_9 ? 4'h9 : _reqChosen_T_4; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_6 = reqIdleBits_8 ? 4'h8 : _reqChosen_T_5; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_7 = reqIdleBits_7 ? 4'h7 : _reqChosen_T_6; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_8 = reqIdleBits_6 ? 4'h6 : _reqChosen_T_7; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_9 = reqIdleBits_5 ? 4'h5 : _reqChosen_T_8; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_10 = reqIdleBits_4 ? 4'h4 : _reqChosen_T_9; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_11 = reqIdleBits_3 ? 4'h3 : _reqChosen_T_10; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_12 = reqIdleBits_2 ? 4'h2 : _reqChosen_T_11; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_13 = reqIdleBits_1 ? 4'h1 : _reqChosen_T_12; // @[Mux.scala 47:70]
  wire [3:0] reqChosen = reqIdleBits_0 ? 4'h0 : _reqChosen_T_13; // @[Mux.scala 47:70]
  reg [15:0] req_cache_0_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_1_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_2_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_3_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_4_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_5_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_6_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_7_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_8_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_9_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_10_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_11_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_12_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_13_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_14_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_15_memoryLength; // @[CScratchpad.scala 114:30]
  reg [33:0] totalTx_memoryAddress; // @[CScratchpad.scala 124:28]
  reg [33:0] totalTx_memoryLength; // @[CScratchpad.scala 124:28]
  wire  isBelowLimit = totalTx_memoryLength <= 34'h40; // @[CScratchpad.scala 149:47]
  wire [1:0] txEmitLengthLg_hi = totalTx_memoryLength[33:32]; // @[OneHot.scala 30:18]
  wire  _txEmitLengthLg_T = |txEmitLengthLg_hi; // @[OneHot.scala 32:14]
  wire [31:0] txEmitLengthLg_lo = totalTx_memoryLength[31:0]; // @[OneHot.scala 31:18]
  wire [31:0] _GEN_569 = {{30'd0}, txEmitLengthLg_hi}; // @[OneHot.scala 32:28]
  wire [31:0] _txEmitLengthLg_T_1 = _GEN_569 | txEmitLengthLg_lo; // @[OneHot.scala 32:28]
  wire [15:0] txEmitLengthLg_hi_1 = _txEmitLengthLg_T_1[31:16]; // @[OneHot.scala 30:18]
  wire  _txEmitLengthLg_T_2 = |txEmitLengthLg_hi_1; // @[OneHot.scala 32:14]
  wire [15:0] txEmitLengthLg_lo_1 = _txEmitLengthLg_T_1[15:0]; // @[OneHot.scala 31:18]
  wire [15:0] _txEmitLengthLg_T_3 = txEmitLengthLg_hi_1 | txEmitLengthLg_lo_1; // @[OneHot.scala 32:28]
  wire [7:0] txEmitLengthLg_hi_2 = _txEmitLengthLg_T_3[15:8]; // @[OneHot.scala 30:18]
  wire  _txEmitLengthLg_T_4 = |txEmitLengthLg_hi_2; // @[OneHot.scala 32:14]
  wire [7:0] txEmitLengthLg_lo_2 = _txEmitLengthLg_T_3[7:0]; // @[OneHot.scala 31:18]
  wire [7:0] _txEmitLengthLg_T_5 = txEmitLengthLg_hi_2 | txEmitLengthLg_lo_2; // @[OneHot.scala 32:28]
  wire [3:0] txEmitLengthLg_hi_3 = _txEmitLengthLg_T_5[7:4]; // @[OneHot.scala 30:18]
  wire  _txEmitLengthLg_T_6 = |txEmitLengthLg_hi_3; // @[OneHot.scala 32:14]
  wire [3:0] txEmitLengthLg_lo_3 = _txEmitLengthLg_T_5[3:0]; // @[OneHot.scala 31:18]
  wire [3:0] _txEmitLengthLg_T_7 = txEmitLengthLg_hi_3 | txEmitLengthLg_lo_3; // @[OneHot.scala 32:28]
  wire [1:0] txEmitLengthLg_hi_4 = _txEmitLengthLg_T_7[3:2]; // @[OneHot.scala 30:18]
  wire  _txEmitLengthLg_T_8 = |txEmitLengthLg_hi_4; // @[OneHot.scala 32:14]
  wire [1:0] txEmitLengthLg_lo_4 = _txEmitLengthLg_T_7[1:0]; // @[OneHot.scala 31:18]
  wire [1:0] _txEmitLengthLg_T_9 = txEmitLengthLg_hi_4 | txEmitLengthLg_lo_4; // @[OneHot.scala 32:28]
  wire [5:0] _txEmitLengthLg_T_15 = {_txEmitLengthLg_T,_txEmitLengthLg_T_2,_txEmitLengthLg_T_4,_txEmitLengthLg_T_6,
    _txEmitLengthLg_T_8,_txEmitLengthLg_T_9[1]}; // @[Cat.scala 33:92]
  wire [5:0] _txEmitLengthLg_T_16 = isBelowLimit ? _txEmitLengthLg_T_15 : 6'h6; // @[CScratchpad.scala 150:28]
  wire [5:0] _GEN_111 = 2'h1 == mem_tx_state ? _txEmitLengthLg_T_16 : 6'h0; // @[CScratchpad.scala 131:18 138:24 150:22]
  wire [5:0] _GEN_169 = 2'h0 == mem_tx_state ? 6'h0 : _GEN_111; // @[CScratchpad.scala 131:18 138:24]
  wire [3:0] txEmitLengthLg = _GEN_169[3:0]; // @[CScratchpad.scala 130:36]
  wire [5:0] _x1_a_bits_a_mask_sizeOH_T = {{2'd0}, txEmitLengthLg}; // @[Misc.scala 201:34]
  wire [2:0] x1_a_bits_a_mask_sizeOH_shiftAmount = _x1_a_bits_a_mask_sizeOH_T[2:0]; // @[OneHot.scala 63:49]
  wire [7:0] _x1_a_bits_a_mask_sizeOH_T_1 = 8'h1 << x1_a_bits_a_mask_sizeOH_shiftAmount; // @[OneHot.scala 64:12]
  wire [5:0] x1_a_bits_a_mask_sizeOH = _x1_a_bits_a_mask_sizeOH_T_1[5:0] | 6'h1; // @[Misc.scala 201:81]
  wire  _x1_a_bits_a_mask_T = txEmitLengthLg >= 4'h6; // @[Misc.scala 205:21]
  wire  x1_a_bits_a_mask_size = x1_a_bits_a_mask_sizeOH[5]; // @[Misc.scala 208:26]
  wire  x1_a_bits_a_mask_bit = totalTx_memoryAddress[5]; // @[Misc.scala 209:26]
  wire  x1_a_bits_a_mask_nbit = ~x1_a_bits_a_mask_bit; // @[Misc.scala 210:20]
  wire  x1_a_bits_a_mask_acc = _x1_a_bits_a_mask_T | x1_a_bits_a_mask_size & x1_a_bits_a_mask_nbit; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_acc_1 = _x1_a_bits_a_mask_T | x1_a_bits_a_mask_size & x1_a_bits_a_mask_bit; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_size_1 = x1_a_bits_a_mask_sizeOH[4]; // @[Misc.scala 208:26]
  wire  x1_a_bits_a_mask_bit_1 = totalTx_memoryAddress[4]; // @[Misc.scala 209:26]
  wire  x1_a_bits_a_mask_nbit_1 = ~x1_a_bits_a_mask_bit_1; // @[Misc.scala 210:20]
  wire  x1_a_bits_a_mask_eq_2 = x1_a_bits_a_mask_nbit & x1_a_bits_a_mask_nbit_1; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_2 = x1_a_bits_a_mask_acc | x1_a_bits_a_mask_size_1 & x1_a_bits_a_mask_eq_2; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_3 = x1_a_bits_a_mask_nbit & x1_a_bits_a_mask_bit_1; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_3 = x1_a_bits_a_mask_acc | x1_a_bits_a_mask_size_1 & x1_a_bits_a_mask_eq_3; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_4 = x1_a_bits_a_mask_bit & x1_a_bits_a_mask_nbit_1; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_4 = x1_a_bits_a_mask_acc_1 | x1_a_bits_a_mask_size_1 & x1_a_bits_a_mask_eq_4; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_5 = x1_a_bits_a_mask_bit & x1_a_bits_a_mask_bit_1; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_5 = x1_a_bits_a_mask_acc_1 | x1_a_bits_a_mask_size_1 & x1_a_bits_a_mask_eq_5; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_size_2 = x1_a_bits_a_mask_sizeOH[3]; // @[Misc.scala 208:26]
  wire  x1_a_bits_a_mask_bit_2 = totalTx_memoryAddress[3]; // @[Misc.scala 209:26]
  wire  x1_a_bits_a_mask_nbit_2 = ~x1_a_bits_a_mask_bit_2; // @[Misc.scala 210:20]
  wire  x1_a_bits_a_mask_eq_6 = x1_a_bits_a_mask_eq_2 & x1_a_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_6 = x1_a_bits_a_mask_acc_2 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_6; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_7 = x1_a_bits_a_mask_eq_2 & x1_a_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_7 = x1_a_bits_a_mask_acc_2 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_7; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_8 = x1_a_bits_a_mask_eq_3 & x1_a_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_8 = x1_a_bits_a_mask_acc_3 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_8; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_9 = x1_a_bits_a_mask_eq_3 & x1_a_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_9 = x1_a_bits_a_mask_acc_3 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_9; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_10 = x1_a_bits_a_mask_eq_4 & x1_a_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_10 = x1_a_bits_a_mask_acc_4 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_10; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_11 = x1_a_bits_a_mask_eq_4 & x1_a_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_11 = x1_a_bits_a_mask_acc_4 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_11; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_12 = x1_a_bits_a_mask_eq_5 & x1_a_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_12 = x1_a_bits_a_mask_acc_5 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_12; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_13 = x1_a_bits_a_mask_eq_5 & x1_a_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_13 = x1_a_bits_a_mask_acc_5 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_13; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_size_3 = x1_a_bits_a_mask_sizeOH[2]; // @[Misc.scala 208:26]
  wire  x1_a_bits_a_mask_bit_3 = totalTx_memoryAddress[2]; // @[Misc.scala 209:26]
  wire  x1_a_bits_a_mask_nbit_3 = ~x1_a_bits_a_mask_bit_3; // @[Misc.scala 210:20]
  wire  x1_a_bits_a_mask_eq_14 = x1_a_bits_a_mask_eq_6 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_14 = x1_a_bits_a_mask_acc_6 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_14; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_15 = x1_a_bits_a_mask_eq_6 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_15 = x1_a_bits_a_mask_acc_6 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_15; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_16 = x1_a_bits_a_mask_eq_7 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_16 = x1_a_bits_a_mask_acc_7 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_16; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_17 = x1_a_bits_a_mask_eq_7 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_17 = x1_a_bits_a_mask_acc_7 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_17; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_18 = x1_a_bits_a_mask_eq_8 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_18 = x1_a_bits_a_mask_acc_8 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_18; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_19 = x1_a_bits_a_mask_eq_8 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_19 = x1_a_bits_a_mask_acc_8 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_19; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_20 = x1_a_bits_a_mask_eq_9 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_20 = x1_a_bits_a_mask_acc_9 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_20; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_21 = x1_a_bits_a_mask_eq_9 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_21 = x1_a_bits_a_mask_acc_9 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_21; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_22 = x1_a_bits_a_mask_eq_10 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_22 = x1_a_bits_a_mask_acc_10 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_22; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_23 = x1_a_bits_a_mask_eq_10 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_23 = x1_a_bits_a_mask_acc_10 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_23; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_24 = x1_a_bits_a_mask_eq_11 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_24 = x1_a_bits_a_mask_acc_11 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_24; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_25 = x1_a_bits_a_mask_eq_11 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_25 = x1_a_bits_a_mask_acc_11 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_25; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_26 = x1_a_bits_a_mask_eq_12 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_26 = x1_a_bits_a_mask_acc_12 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_26; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_27 = x1_a_bits_a_mask_eq_12 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_27 = x1_a_bits_a_mask_acc_12 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_27; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_28 = x1_a_bits_a_mask_eq_13 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_28 = x1_a_bits_a_mask_acc_13 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_28; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_29 = x1_a_bits_a_mask_eq_13 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_29 = x1_a_bits_a_mask_acc_13 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_29; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_size_4 = x1_a_bits_a_mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  x1_a_bits_a_mask_bit_4 = totalTx_memoryAddress[1]; // @[Misc.scala 209:26]
  wire  x1_a_bits_a_mask_nbit_4 = ~x1_a_bits_a_mask_bit_4; // @[Misc.scala 210:20]
  wire  x1_a_bits_a_mask_eq_30 = x1_a_bits_a_mask_eq_14 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_30 = x1_a_bits_a_mask_acc_14 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_30; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_31 = x1_a_bits_a_mask_eq_14 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_31 = x1_a_bits_a_mask_acc_14 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_31; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_32 = x1_a_bits_a_mask_eq_15 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_32 = x1_a_bits_a_mask_acc_15 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_32; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_33 = x1_a_bits_a_mask_eq_15 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_33 = x1_a_bits_a_mask_acc_15 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_33; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_34 = x1_a_bits_a_mask_eq_16 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_34 = x1_a_bits_a_mask_acc_16 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_34; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_35 = x1_a_bits_a_mask_eq_16 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_35 = x1_a_bits_a_mask_acc_16 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_35; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_36 = x1_a_bits_a_mask_eq_17 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_36 = x1_a_bits_a_mask_acc_17 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_36; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_37 = x1_a_bits_a_mask_eq_17 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_37 = x1_a_bits_a_mask_acc_17 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_37; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_38 = x1_a_bits_a_mask_eq_18 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_38 = x1_a_bits_a_mask_acc_18 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_38; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_39 = x1_a_bits_a_mask_eq_18 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_39 = x1_a_bits_a_mask_acc_18 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_39; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_40 = x1_a_bits_a_mask_eq_19 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_40 = x1_a_bits_a_mask_acc_19 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_40; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_41 = x1_a_bits_a_mask_eq_19 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_41 = x1_a_bits_a_mask_acc_19 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_41; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_42 = x1_a_bits_a_mask_eq_20 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_42 = x1_a_bits_a_mask_acc_20 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_42; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_43 = x1_a_bits_a_mask_eq_20 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_43 = x1_a_bits_a_mask_acc_20 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_43; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_44 = x1_a_bits_a_mask_eq_21 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_44 = x1_a_bits_a_mask_acc_21 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_44; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_45 = x1_a_bits_a_mask_eq_21 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_45 = x1_a_bits_a_mask_acc_21 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_45; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_46 = x1_a_bits_a_mask_eq_22 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_46 = x1_a_bits_a_mask_acc_22 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_46; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_47 = x1_a_bits_a_mask_eq_22 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_47 = x1_a_bits_a_mask_acc_22 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_47; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_48 = x1_a_bits_a_mask_eq_23 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_48 = x1_a_bits_a_mask_acc_23 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_48; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_49 = x1_a_bits_a_mask_eq_23 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_49 = x1_a_bits_a_mask_acc_23 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_49; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_50 = x1_a_bits_a_mask_eq_24 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_50 = x1_a_bits_a_mask_acc_24 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_50; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_51 = x1_a_bits_a_mask_eq_24 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_51 = x1_a_bits_a_mask_acc_24 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_51; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_52 = x1_a_bits_a_mask_eq_25 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_52 = x1_a_bits_a_mask_acc_25 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_52; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_53 = x1_a_bits_a_mask_eq_25 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_53 = x1_a_bits_a_mask_acc_25 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_53; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_54 = x1_a_bits_a_mask_eq_26 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_54 = x1_a_bits_a_mask_acc_26 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_54; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_55 = x1_a_bits_a_mask_eq_26 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_55 = x1_a_bits_a_mask_acc_26 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_55; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_56 = x1_a_bits_a_mask_eq_27 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_56 = x1_a_bits_a_mask_acc_27 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_56; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_57 = x1_a_bits_a_mask_eq_27 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_57 = x1_a_bits_a_mask_acc_27 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_57; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_58 = x1_a_bits_a_mask_eq_28 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_58 = x1_a_bits_a_mask_acc_28 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_58; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_59 = x1_a_bits_a_mask_eq_28 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_59 = x1_a_bits_a_mask_acc_28 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_59; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_60 = x1_a_bits_a_mask_eq_29 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_60 = x1_a_bits_a_mask_acc_29 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_60; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_61 = x1_a_bits_a_mask_eq_29 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_61 = x1_a_bits_a_mask_acc_29 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_61; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_size_5 = x1_a_bits_a_mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  x1_a_bits_a_mask_bit_5 = totalTx_memoryAddress[0]; // @[Misc.scala 209:26]
  wire  x1_a_bits_a_mask_nbit_5 = ~x1_a_bits_a_mask_bit_5; // @[Misc.scala 210:20]
  wire  x1_a_bits_a_mask_eq_62 = x1_a_bits_a_mask_eq_30 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_62 = x1_a_bits_a_mask_acc_30 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_62; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_63 = x1_a_bits_a_mask_eq_30 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_63 = x1_a_bits_a_mask_acc_30 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_63; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_64 = x1_a_bits_a_mask_eq_31 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_64 = x1_a_bits_a_mask_acc_31 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_64; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_65 = x1_a_bits_a_mask_eq_31 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_65 = x1_a_bits_a_mask_acc_31 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_65; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_66 = x1_a_bits_a_mask_eq_32 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_66 = x1_a_bits_a_mask_acc_32 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_66; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_67 = x1_a_bits_a_mask_eq_32 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_67 = x1_a_bits_a_mask_acc_32 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_67; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_68 = x1_a_bits_a_mask_eq_33 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_68 = x1_a_bits_a_mask_acc_33 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_68; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_69 = x1_a_bits_a_mask_eq_33 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_69 = x1_a_bits_a_mask_acc_33 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_69; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_70 = x1_a_bits_a_mask_eq_34 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_70 = x1_a_bits_a_mask_acc_34 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_70; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_71 = x1_a_bits_a_mask_eq_34 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_71 = x1_a_bits_a_mask_acc_34 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_71; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_72 = x1_a_bits_a_mask_eq_35 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_72 = x1_a_bits_a_mask_acc_35 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_72; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_73 = x1_a_bits_a_mask_eq_35 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_73 = x1_a_bits_a_mask_acc_35 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_73; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_74 = x1_a_bits_a_mask_eq_36 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_74 = x1_a_bits_a_mask_acc_36 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_74; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_75 = x1_a_bits_a_mask_eq_36 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_75 = x1_a_bits_a_mask_acc_36 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_75; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_76 = x1_a_bits_a_mask_eq_37 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_76 = x1_a_bits_a_mask_acc_37 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_76; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_77 = x1_a_bits_a_mask_eq_37 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_77 = x1_a_bits_a_mask_acc_37 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_77; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_78 = x1_a_bits_a_mask_eq_38 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_78 = x1_a_bits_a_mask_acc_38 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_78; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_79 = x1_a_bits_a_mask_eq_38 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_79 = x1_a_bits_a_mask_acc_38 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_79; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_80 = x1_a_bits_a_mask_eq_39 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_80 = x1_a_bits_a_mask_acc_39 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_80; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_81 = x1_a_bits_a_mask_eq_39 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_81 = x1_a_bits_a_mask_acc_39 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_81; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_82 = x1_a_bits_a_mask_eq_40 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_82 = x1_a_bits_a_mask_acc_40 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_82; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_83 = x1_a_bits_a_mask_eq_40 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_83 = x1_a_bits_a_mask_acc_40 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_83; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_84 = x1_a_bits_a_mask_eq_41 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_84 = x1_a_bits_a_mask_acc_41 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_84; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_85 = x1_a_bits_a_mask_eq_41 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_85 = x1_a_bits_a_mask_acc_41 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_85; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_86 = x1_a_bits_a_mask_eq_42 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_86 = x1_a_bits_a_mask_acc_42 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_86; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_87 = x1_a_bits_a_mask_eq_42 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_87 = x1_a_bits_a_mask_acc_42 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_87; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_88 = x1_a_bits_a_mask_eq_43 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_88 = x1_a_bits_a_mask_acc_43 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_88; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_89 = x1_a_bits_a_mask_eq_43 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_89 = x1_a_bits_a_mask_acc_43 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_89; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_90 = x1_a_bits_a_mask_eq_44 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_90 = x1_a_bits_a_mask_acc_44 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_90; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_91 = x1_a_bits_a_mask_eq_44 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_91 = x1_a_bits_a_mask_acc_44 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_91; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_92 = x1_a_bits_a_mask_eq_45 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_92 = x1_a_bits_a_mask_acc_45 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_92; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_93 = x1_a_bits_a_mask_eq_45 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_93 = x1_a_bits_a_mask_acc_45 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_93; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_94 = x1_a_bits_a_mask_eq_46 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_94 = x1_a_bits_a_mask_acc_46 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_94; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_95 = x1_a_bits_a_mask_eq_46 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_95 = x1_a_bits_a_mask_acc_46 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_95; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_96 = x1_a_bits_a_mask_eq_47 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_96 = x1_a_bits_a_mask_acc_47 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_96; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_97 = x1_a_bits_a_mask_eq_47 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_97 = x1_a_bits_a_mask_acc_47 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_97; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_98 = x1_a_bits_a_mask_eq_48 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_98 = x1_a_bits_a_mask_acc_48 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_98; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_99 = x1_a_bits_a_mask_eq_48 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_99 = x1_a_bits_a_mask_acc_48 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_99; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_100 = x1_a_bits_a_mask_eq_49 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_100 = x1_a_bits_a_mask_acc_49 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_100; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_101 = x1_a_bits_a_mask_eq_49 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_101 = x1_a_bits_a_mask_acc_49 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_101; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_102 = x1_a_bits_a_mask_eq_50 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_102 = x1_a_bits_a_mask_acc_50 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_102; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_103 = x1_a_bits_a_mask_eq_50 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_103 = x1_a_bits_a_mask_acc_50 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_103; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_104 = x1_a_bits_a_mask_eq_51 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_104 = x1_a_bits_a_mask_acc_51 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_104; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_105 = x1_a_bits_a_mask_eq_51 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_105 = x1_a_bits_a_mask_acc_51 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_105; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_106 = x1_a_bits_a_mask_eq_52 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_106 = x1_a_bits_a_mask_acc_52 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_106; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_107 = x1_a_bits_a_mask_eq_52 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_107 = x1_a_bits_a_mask_acc_52 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_107; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_108 = x1_a_bits_a_mask_eq_53 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_108 = x1_a_bits_a_mask_acc_53 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_108; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_109 = x1_a_bits_a_mask_eq_53 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_109 = x1_a_bits_a_mask_acc_53 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_109; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_110 = x1_a_bits_a_mask_eq_54 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_110 = x1_a_bits_a_mask_acc_54 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_110; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_111 = x1_a_bits_a_mask_eq_54 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_111 = x1_a_bits_a_mask_acc_54 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_111; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_112 = x1_a_bits_a_mask_eq_55 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_112 = x1_a_bits_a_mask_acc_55 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_112; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_113 = x1_a_bits_a_mask_eq_55 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_113 = x1_a_bits_a_mask_acc_55 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_113; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_114 = x1_a_bits_a_mask_eq_56 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_114 = x1_a_bits_a_mask_acc_56 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_114; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_115 = x1_a_bits_a_mask_eq_56 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_115 = x1_a_bits_a_mask_acc_56 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_115; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_116 = x1_a_bits_a_mask_eq_57 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_116 = x1_a_bits_a_mask_acc_57 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_116; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_117 = x1_a_bits_a_mask_eq_57 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_117 = x1_a_bits_a_mask_acc_57 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_117; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_118 = x1_a_bits_a_mask_eq_58 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_118 = x1_a_bits_a_mask_acc_58 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_118; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_119 = x1_a_bits_a_mask_eq_58 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_119 = x1_a_bits_a_mask_acc_58 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_119; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_120 = x1_a_bits_a_mask_eq_59 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_120 = x1_a_bits_a_mask_acc_59 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_120; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_121 = x1_a_bits_a_mask_eq_59 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_121 = x1_a_bits_a_mask_acc_59 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_121; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_122 = x1_a_bits_a_mask_eq_60 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_122 = x1_a_bits_a_mask_acc_60 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_122; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_123 = x1_a_bits_a_mask_eq_60 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_123 = x1_a_bits_a_mask_acc_60 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_123; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_124 = x1_a_bits_a_mask_eq_61 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_124 = x1_a_bits_a_mask_acc_61 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_124; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_125 = x1_a_bits_a_mask_eq_61 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_125 = x1_a_bits_a_mask_acc_61 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_125; // @[Misc.scala 214:29]
  wire [7:0] x1_a_bits_a_mask_lo_lo_lo = {x1_a_bits_a_mask_acc_69,x1_a_bits_a_mask_acc_68,x1_a_bits_a_mask_acc_67,
    x1_a_bits_a_mask_acc_66,x1_a_bits_a_mask_acc_65,x1_a_bits_a_mask_acc_64,x1_a_bits_a_mask_acc_63,
    x1_a_bits_a_mask_acc_62}; // @[Cat.scala 33:92]
  wire [15:0] x1_a_bits_a_mask_lo_lo = {x1_a_bits_a_mask_acc_77,x1_a_bits_a_mask_acc_76,x1_a_bits_a_mask_acc_75,
    x1_a_bits_a_mask_acc_74,x1_a_bits_a_mask_acc_73,x1_a_bits_a_mask_acc_72,x1_a_bits_a_mask_acc_71,
    x1_a_bits_a_mask_acc_70,x1_a_bits_a_mask_lo_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] x1_a_bits_a_mask_lo_hi_lo = {x1_a_bits_a_mask_acc_85,x1_a_bits_a_mask_acc_84,x1_a_bits_a_mask_acc_83,
    x1_a_bits_a_mask_acc_82,x1_a_bits_a_mask_acc_81,x1_a_bits_a_mask_acc_80,x1_a_bits_a_mask_acc_79,
    x1_a_bits_a_mask_acc_78}; // @[Cat.scala 33:92]
  wire [31:0] x1_a_bits_a_mask_lo = {x1_a_bits_a_mask_acc_93,x1_a_bits_a_mask_acc_92,x1_a_bits_a_mask_acc_91,
    x1_a_bits_a_mask_acc_90,x1_a_bits_a_mask_acc_89,x1_a_bits_a_mask_acc_88,x1_a_bits_a_mask_acc_87,
    x1_a_bits_a_mask_acc_86,x1_a_bits_a_mask_lo_hi_lo,x1_a_bits_a_mask_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] x1_a_bits_a_mask_hi_lo_lo = {x1_a_bits_a_mask_acc_101,x1_a_bits_a_mask_acc_100,x1_a_bits_a_mask_acc_99,
    x1_a_bits_a_mask_acc_98,x1_a_bits_a_mask_acc_97,x1_a_bits_a_mask_acc_96,x1_a_bits_a_mask_acc_95,
    x1_a_bits_a_mask_acc_94}; // @[Cat.scala 33:92]
  wire [15:0] x1_a_bits_a_mask_hi_lo = {x1_a_bits_a_mask_acc_109,x1_a_bits_a_mask_acc_108,x1_a_bits_a_mask_acc_107,
    x1_a_bits_a_mask_acc_106,x1_a_bits_a_mask_acc_105,x1_a_bits_a_mask_acc_104,x1_a_bits_a_mask_acc_103,
    x1_a_bits_a_mask_acc_102,x1_a_bits_a_mask_hi_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] x1_a_bits_a_mask_hi_hi_lo = {x1_a_bits_a_mask_acc_117,x1_a_bits_a_mask_acc_116,x1_a_bits_a_mask_acc_115,
    x1_a_bits_a_mask_acc_114,x1_a_bits_a_mask_acc_113,x1_a_bits_a_mask_acc_112,x1_a_bits_a_mask_acc_111,
    x1_a_bits_a_mask_acc_110}; // @[Cat.scala 33:92]
  wire [31:0] x1_a_bits_a_mask_hi = {x1_a_bits_a_mask_acc_125,x1_a_bits_a_mask_acc_124,x1_a_bits_a_mask_acc_123,
    x1_a_bits_a_mask_acc_122,x1_a_bits_a_mask_acc_121,x1_a_bits_a_mask_acc_120,x1_a_bits_a_mask_acc_119,
    x1_a_bits_a_mask_acc_118,x1_a_bits_a_mask_hi_hi_lo,x1_a_bits_a_mask_hi_lo}; // @[Cat.scala 33:92]
  wire  _GEN_112 = 2'h1 == mem_tx_state ? reqAvailable : mem_tx_state == 2'h1; // @[CScratchpad.scala 136:19 138:24 151:23]
  wire  mem_out_a_valid = 2'h0 == mem_tx_state ? mem_tx_state == 2'h1 : _GEN_112; // @[CScratchpad.scala 136:19 138:24]
  wire  _T_13 = auto_mem_out_a_ready & mem_out_a_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_8 = 4'h0 == reqChosen ? 1'h0 : reqIdleBits_0; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_9 = 4'h1 == reqChosen ? 1'h0 : reqIdleBits_1; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_10 = 4'h2 == reqChosen ? 1'h0 : reqIdleBits_2; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_11 = 4'h3 == reqChosen ? 1'h0 : reqIdleBits_3; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_12 = 4'h4 == reqChosen ? 1'h0 : reqIdleBits_4; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_13 = 4'h5 == reqChosen ? 1'h0 : reqIdleBits_5; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_14 = 4'h6 == reqChosen ? 1'h0 : reqIdleBits_6; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_15 = 4'h7 == reqChosen ? 1'h0 : reqIdleBits_7; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_16 = 4'h8 == reqChosen ? 1'h0 : reqIdleBits_8; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_17 = 4'h9 == reqChosen ? 1'h0 : reqIdleBits_9; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_18 = 4'ha == reqChosen ? 1'h0 : reqIdleBits_10; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_19 = 4'hb == reqChosen ? 1'h0 : reqIdleBits_11; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_20 = 4'hc == reqChosen ? 1'h0 : reqIdleBits_12; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_21 = 4'hd == reqChosen ? 1'h0 : reqIdleBits_13; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_22 = 4'he == reqChosen ? 1'h0 : reqIdleBits_14; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_23 = 4'hf == reqChosen ? 1'h0 : reqIdleBits_15; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire [33:0] _req_cache_memoryLength_T = isBelowLimit ? totalTx_memoryLength : 34'h40; // @[CScratchpad.scala 155:49]
  wire [15:0] _GEN_40 = 4'h0 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_0_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_41 = 4'h1 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_1_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_42 = 4'h2 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_2_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_43 = 4'h3 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_3_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_44 = 4'h4 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_4_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_45 = 4'h5 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_5_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_46 = 4'h6 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_6_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_47 = 4'h7 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_7_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_48 = 4'h8 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_8_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_49 = 4'h9 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_9_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_50 = 4'ha == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_10_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_51 = 4'hb == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_11_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_52 = 4'hc == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_12_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_53 = 4'hd == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_13_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_54 = 4'he == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_14_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_55 = 4'hf == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_15_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [33:0] _totalTx_memoryLength_T_1 = totalTx_memoryLength - 34'h40; // @[CScratchpad.scala 156:54]
  wire [33:0] _totalTx_memoryAddress_T_1 = totalTx_memoryAddress + 34'h40; // @[CScratchpad.scala 158:56]
  wire [1:0] _GEN_56 = isBelowLimit ? 2'h2 : mem_tx_state; // @[CScratchpad.scala 159:28 160:24 102:37]
  wire  _GEN_57 = _T_13 ? _GEN_8 : reqIdleBits_0; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_58 = _T_13 ? _GEN_9 : reqIdleBits_1; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_59 = _T_13 ? _GEN_10 : reqIdleBits_2; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_60 = _T_13 ? _GEN_11 : reqIdleBits_3; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_61 = _T_13 ? _GEN_12 : reqIdleBits_4; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_62 = _T_13 ? _GEN_13 : reqIdleBits_5; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_63 = _T_13 ? _GEN_14 : reqIdleBits_6; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_64 = _T_13 ? _GEN_15 : reqIdleBits_7; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_65 = _T_13 ? _GEN_16 : reqIdleBits_8; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_66 = _T_13 ? _GEN_17 : reqIdleBits_9; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_67 = _T_13 ? _GEN_18 : reqIdleBits_10; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_68 = _T_13 ? _GEN_19 : reqIdleBits_11; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_69 = _T_13 ? _GEN_20 : reqIdleBits_12; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_70 = _T_13 ? _GEN_21 : reqIdleBits_13; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_71 = _T_13 ? _GEN_22 : reqIdleBits_14; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_72 = _T_13 ? _GEN_23 : reqIdleBits_15; // @[CScratchpad.scala 152:28 110:36]
  wire [15:0] _GEN_89 = _T_13 ? _GEN_40 : req_cache_0_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_90 = _T_13 ? _GEN_41 : req_cache_1_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_91 = _T_13 ? _GEN_42 : req_cache_2_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_92 = _T_13 ? _GEN_43 : req_cache_3_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_93 = _T_13 ? _GEN_44 : req_cache_4_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_94 = _T_13 ? _GEN_45 : req_cache_5_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_95 = _T_13 ? _GEN_46 : req_cache_6_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_96 = _T_13 ? _GEN_47 : req_cache_7_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_97 = _T_13 ? _GEN_48 : req_cache_8_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_98 = _T_13 ? _GEN_49 : req_cache_9_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_99 = _T_13 ? _GEN_50 : req_cache_10_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_100 = _T_13 ? _GEN_51 : req_cache_11_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_101 = _T_13 ? _GEN_52 : req_cache_12_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_102 = _T_13 ? _GEN_53 : req_cache_13_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_103 = _T_13 ? _GEN_54 : req_cache_14_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_104 = _T_13 ? _GEN_55 : req_cache_15_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [1:0] _GEN_109 = reqIdleBits_0 & reqIdleBits_1 & reqIdleBits_2 & reqIdleBits_3 & reqIdleBits_4 & reqIdleBits_5 &
    reqIdleBits_6 & reqIdleBits_7 & reqIdleBits_8 & reqIdleBits_9 & reqIdleBits_10 & reqIdleBits_11 & reqIdleBits_12 &
    reqIdleBits_13 & reqIdleBits_14 & reqIdleBits_15 ? 2'h0 : mem_tx_state; // @[CScratchpad.scala 166:40 167:22 102:37]
  wire  _GEN_113 = 2'h1 == mem_tx_state ? _GEN_57 : reqIdleBits_0; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_114 = 2'h1 == mem_tx_state ? _GEN_58 : reqIdleBits_1; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_115 = 2'h1 == mem_tx_state ? _GEN_59 : reqIdleBits_2; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_116 = 2'h1 == mem_tx_state ? _GEN_60 : reqIdleBits_3; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_117 = 2'h1 == mem_tx_state ? _GEN_61 : reqIdleBits_4; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_118 = 2'h1 == mem_tx_state ? _GEN_62 : reqIdleBits_5; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_119 = 2'h1 == mem_tx_state ? _GEN_63 : reqIdleBits_6; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_120 = 2'h1 == mem_tx_state ? _GEN_64 : reqIdleBits_7; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_121 = 2'h1 == mem_tx_state ? _GEN_65 : reqIdleBits_8; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_122 = 2'h1 == mem_tx_state ? _GEN_66 : reqIdleBits_9; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_123 = 2'h1 == mem_tx_state ? _GEN_67 : reqIdleBits_10; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_124 = 2'h1 == mem_tx_state ? _GEN_68 : reqIdleBits_11; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_125 = 2'h1 == mem_tx_state ? _GEN_69 : reqIdleBits_12; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_126 = 2'h1 == mem_tx_state ? _GEN_70 : reqIdleBits_13; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_127 = 2'h1 == mem_tx_state ? _GEN_71 : reqIdleBits_14; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_128 = 2'h1 == mem_tx_state ? _GEN_72 : reqIdleBits_15; // @[CScratchpad.scala 138:24 110:36]
  wire [15:0] _GEN_145 = 2'h1 == mem_tx_state ? _GEN_89 : req_cache_0_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_146 = 2'h1 == mem_tx_state ? _GEN_90 : req_cache_1_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_147 = 2'h1 == mem_tx_state ? _GEN_91 : req_cache_2_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_148 = 2'h1 == mem_tx_state ? _GEN_92 : req_cache_3_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_149 = 2'h1 == mem_tx_state ? _GEN_93 : req_cache_4_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_150 = 2'h1 == mem_tx_state ? _GEN_94 : req_cache_5_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_151 = 2'h1 == mem_tx_state ? _GEN_95 : req_cache_6_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_152 = 2'h1 == mem_tx_state ? _GEN_96 : req_cache_7_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_153 = 2'h1 == mem_tx_state ? _GEN_97 : req_cache_8_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_154 = 2'h1 == mem_tx_state ? _GEN_98 : req_cache_9_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_155 = 2'h1 == mem_tx_state ? _GEN_99 : req_cache_10_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_156 = 2'h1 == mem_tx_state ? _GEN_100 : req_cache_11_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_157 = 2'h1 == mem_tx_state ? _GEN_101 : req_cache_12_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_158 = 2'h1 == mem_tx_state ? _GEN_102 : req_cache_13_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_159 = 2'h1 == mem_tx_state ? _GEN_103 : req_cache_14_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_160 = 2'h1 == mem_tx_state ? _GEN_104 : req_cache_15_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire  _GEN_171 = 2'h0 == mem_tx_state ? reqIdleBits_0 : _GEN_113; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_172 = 2'h0 == mem_tx_state ? reqIdleBits_1 : _GEN_114; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_173 = 2'h0 == mem_tx_state ? reqIdleBits_2 : _GEN_115; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_174 = 2'h0 == mem_tx_state ? reqIdleBits_3 : _GEN_116; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_175 = 2'h0 == mem_tx_state ? reqIdleBits_4 : _GEN_117; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_176 = 2'h0 == mem_tx_state ? reqIdleBits_5 : _GEN_118; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_177 = 2'h0 == mem_tx_state ? reqIdleBits_6 : _GEN_119; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_178 = 2'h0 == mem_tx_state ? reqIdleBits_7 : _GEN_120; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_179 = 2'h0 == mem_tx_state ? reqIdleBits_8 : _GEN_121; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_180 = 2'h0 == mem_tx_state ? reqIdleBits_9 : _GEN_122; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_181 = 2'h0 == mem_tx_state ? reqIdleBits_10 : _GEN_123; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_182 = 2'h0 == mem_tx_state ? reqIdleBits_11 : _GEN_124; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_183 = 2'h0 == mem_tx_state ? reqIdleBits_12 : _GEN_125; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_184 = 2'h0 == mem_tx_state ? reqIdleBits_13 : _GEN_126; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_185 = 2'h0 == mem_tx_state ? reqIdleBits_14 : _GEN_127; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_186 = 2'h0 == mem_tx_state ? reqIdleBits_15 : _GEN_128; // @[CScratchpad.scala 138:24 110:36]
  wire [15:0] _GEN_203 = 2'h0 == mem_tx_state ? req_cache_0_memoryLength : _GEN_145; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_204 = 2'h0 == mem_tx_state ? req_cache_1_memoryLength : _GEN_146; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_205 = 2'h0 == mem_tx_state ? req_cache_2_memoryLength : _GEN_147; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_206 = 2'h0 == mem_tx_state ? req_cache_3_memoryLength : _GEN_148; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_207 = 2'h0 == mem_tx_state ? req_cache_4_memoryLength : _GEN_149; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_208 = 2'h0 == mem_tx_state ? req_cache_5_memoryLength : _GEN_150; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_209 = 2'h0 == mem_tx_state ? req_cache_6_memoryLength : _GEN_151; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_210 = 2'h0 == mem_tx_state ? req_cache_7_memoryLength : _GEN_152; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_211 = 2'h0 == mem_tx_state ? req_cache_8_memoryLength : _GEN_153; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_212 = 2'h0 == mem_tx_state ? req_cache_9_memoryLength : _GEN_154; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_213 = 2'h0 == mem_tx_state ? req_cache_10_memoryLength : _GEN_155; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_214 = 2'h0 == mem_tx_state ? req_cache_11_memoryLength : _GEN_156; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_215 = 2'h0 == mem_tx_state ? req_cache_12_memoryLength : _GEN_157; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_216 = 2'h0 == mem_tx_state ? req_cache_13_memoryLength : _GEN_158; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_217 = 2'h0 == mem_tx_state ? req_cache_14_memoryLength : _GEN_159; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_218 = 2'h0 == mem_tx_state ? req_cache_15_memoryLength : _GEN_160; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_220 = 4'h1 == auto_mem_out_d_bits_source ? req_cache_1_memoryLength : req_cache_0_memoryLength; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_221 = 4'h2 == auto_mem_out_d_bits_source ? req_cache_2_memoryLength : _GEN_220; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_222 = 4'h3 == auto_mem_out_d_bits_source ? req_cache_3_memoryLength : _GEN_221; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_223 = 4'h4 == auto_mem_out_d_bits_source ? req_cache_4_memoryLength : _GEN_222; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_224 = 4'h5 == auto_mem_out_d_bits_source ? req_cache_5_memoryLength : _GEN_223; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_225 = 4'h6 == auto_mem_out_d_bits_source ? req_cache_6_memoryLength : _GEN_224; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_226 = 4'h7 == auto_mem_out_d_bits_source ? req_cache_7_memoryLength : _GEN_225; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_227 = 4'h8 == auto_mem_out_d_bits_source ? req_cache_8_memoryLength : _GEN_226; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_228 = 4'h9 == auto_mem_out_d_bits_source ? req_cache_9_memoryLength : _GEN_227; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_229 = 4'ha == auto_mem_out_d_bits_source ? req_cache_10_memoryLength : _GEN_228; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_230 = 4'hb == auto_mem_out_d_bits_source ? req_cache_11_memoryLength : _GEN_229; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_231 = 4'hc == auto_mem_out_d_bits_source ? req_cache_12_memoryLength : _GEN_230; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_232 = 4'hd == auto_mem_out_d_bits_source ? req_cache_13_memoryLength : _GEN_231; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_233 = 4'he == auto_mem_out_d_bits_source ? req_cache_14_memoryLength : _GEN_232; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_234 = 4'hf == auto_mem_out_d_bits_source ? req_cache_15_memoryLength : _GEN_233; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_235 = _GEN_234 >= 16'h40 ? 16'h40 : _GEN_234; // @[CScratchpad.scala 174:55 175:39 177:39]
  wire  mem_out_d_ready = loader_io_cache_block_in_ready; // @[Nodes.scala 1212:84 CScratchpad.scala 180:19]
  wire  _T_36 = mem_out_d_ready & auto_mem_out_d_valid; // @[Decoupled.scala 51:35]
  wire [15:0] _req_cache_memoryLength_T_2 = _GEN_234 - 16'h40; // @[CScratchpad.scala 210:72]
  wire  _GEN_445 = 4'h0 == auto_mem_out_d_bits_source | _GEN_171; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_446 = 4'h1 == auto_mem_out_d_bits_source | _GEN_172; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_447 = 4'h2 == auto_mem_out_d_bits_source | _GEN_173; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_448 = 4'h3 == auto_mem_out_d_bits_source | _GEN_174; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_449 = 4'h4 == auto_mem_out_d_bits_source | _GEN_175; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_450 = 4'h5 == auto_mem_out_d_bits_source | _GEN_176; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_451 = 4'h6 == auto_mem_out_d_bits_source | _GEN_177; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_452 = 4'h7 == auto_mem_out_d_bits_source | _GEN_178; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_453 = 4'h8 == auto_mem_out_d_bits_source | _GEN_179; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_454 = 4'h9 == auto_mem_out_d_bits_source | _GEN_180; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_455 = 4'ha == auto_mem_out_d_bits_source | _GEN_181; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_456 = 4'hb == auto_mem_out_d_bits_source | _GEN_182; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_457 = 4'hc == auto_mem_out_d_bits_source | _GEN_183; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_458 = 4'hd == auto_mem_out_d_bits_source | _GEN_184; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_459 = 4'he == auto_mem_out_d_bits_source | _GEN_185; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_460 = 4'hf == auto_mem_out_d_bits_source | _GEN_186; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_461 = _GEN_234 <= 16'h40 ? _GEN_445 : _GEN_171; // @[CScratchpad.scala 212:57]
  wire  _GEN_462 = _GEN_234 <= 16'h40 ? _GEN_446 : _GEN_172; // @[CScratchpad.scala 212:57]
  wire  _GEN_463 = _GEN_234 <= 16'h40 ? _GEN_447 : _GEN_173; // @[CScratchpad.scala 212:57]
  wire  _GEN_464 = _GEN_234 <= 16'h40 ? _GEN_448 : _GEN_174; // @[CScratchpad.scala 212:57]
  wire  _GEN_465 = _GEN_234 <= 16'h40 ? _GEN_449 : _GEN_175; // @[CScratchpad.scala 212:57]
  wire  _GEN_466 = _GEN_234 <= 16'h40 ? _GEN_450 : _GEN_176; // @[CScratchpad.scala 212:57]
  wire  _GEN_467 = _GEN_234 <= 16'h40 ? _GEN_451 : _GEN_177; // @[CScratchpad.scala 212:57]
  wire  _GEN_468 = _GEN_234 <= 16'h40 ? _GEN_452 : _GEN_178; // @[CScratchpad.scala 212:57]
  wire  _GEN_469 = _GEN_234 <= 16'h40 ? _GEN_453 : _GEN_179; // @[CScratchpad.scala 212:57]
  wire  _GEN_470 = _GEN_234 <= 16'h40 ? _GEN_454 : _GEN_180; // @[CScratchpad.scala 212:57]
  wire  _GEN_471 = _GEN_234 <= 16'h40 ? _GEN_455 : _GEN_181; // @[CScratchpad.scala 212:57]
  wire  _GEN_472 = _GEN_234 <= 16'h40 ? _GEN_456 : _GEN_182; // @[CScratchpad.scala 212:57]
  wire  _GEN_473 = _GEN_234 <= 16'h40 ? _GEN_457 : _GEN_183; // @[CScratchpad.scala 212:57]
  wire  _GEN_474 = _GEN_234 <= 16'h40 ? _GEN_458 : _GEN_184; // @[CScratchpad.scala 212:57]
  wire  _GEN_475 = _GEN_234 <= 16'h40 ? _GEN_459 : _GEN_185; // @[CScratchpad.scala 212:57]
  wire  _GEN_476 = _GEN_234 <= 16'h40 ? _GEN_460 : _GEN_186; // @[CScratchpad.scala 212:57]
  wire  _GEN_494 = _T_36 ? _GEN_461 : _GEN_171; // @[CScratchpad.scala 209:24]
  wire  _GEN_495 = _T_36 ? _GEN_462 : _GEN_172; // @[CScratchpad.scala 209:24]
  wire  _GEN_496 = _T_36 ? _GEN_463 : _GEN_173; // @[CScratchpad.scala 209:24]
  wire  _GEN_497 = _T_36 ? _GEN_464 : _GEN_174; // @[CScratchpad.scala 209:24]
  wire  _GEN_498 = _T_36 ? _GEN_465 : _GEN_175; // @[CScratchpad.scala 209:24]
  wire  _GEN_499 = _T_36 ? _GEN_466 : _GEN_176; // @[CScratchpad.scala 209:24]
  wire  _GEN_500 = _T_36 ? _GEN_467 : _GEN_177; // @[CScratchpad.scala 209:24]
  wire  _GEN_501 = _T_36 ? _GEN_468 : _GEN_178; // @[CScratchpad.scala 209:24]
  wire  _GEN_502 = _T_36 ? _GEN_469 : _GEN_179; // @[CScratchpad.scala 209:24]
  wire  _GEN_503 = _T_36 ? _GEN_470 : _GEN_180; // @[CScratchpad.scala 209:24]
  wire  _GEN_504 = _T_36 ? _GEN_471 : _GEN_181; // @[CScratchpad.scala 209:24]
  wire  _GEN_505 = _T_36 ? _GEN_472 : _GEN_182; // @[CScratchpad.scala 209:24]
  wire  _GEN_506 = _T_36 ? _GEN_473 : _GEN_183; // @[CScratchpad.scala 209:24]
  wire  _GEN_507 = _T_36 ? _GEN_474 : _GEN_184; // @[CScratchpad.scala 209:24]
  wire  _GEN_508 = _T_36 ? _GEN_475 : _GEN_185; // @[CScratchpad.scala 209:24]
  wire  _GEN_509 = _T_36 ? _GEN_476 : _GEN_186; // @[CScratchpad.scala 209:24]
  CScratchpadPackedSubwordLoader_1 loader ( // @[CScratchpad.scala 94:30]
    .clock(loader_clock),
    .reset(loader_reset),
    .io_cache_block_in_ready(loader_io_cache_block_in_ready),
    .io_cache_block_in_valid(loader_io_cache_block_in_valid),
    .io_cache_block_in_bits_len(loader_io_cache_block_in_bits_len),
    .io_sp_write_out_valid(loader_io_sp_write_out_valid)
  );
  assign auto_mem_out_a_valid = 2'h0 == mem_tx_state ? mem_tx_state == 2'h1 : _GEN_112; // @[CScratchpad.scala 136:19 138:24]
  assign auto_mem_out_a_bits_size = txEmitLengthLg[2:0]; // @[Edges.scala 447:17 450:15]
  assign auto_mem_out_a_bits_source = reqIdleBits_0 ? 4'h0 : _reqChosen_T_13; // @[Mux.scala 47:70]
  assign auto_mem_out_a_bits_address = totalTx_memoryAddress; // @[Edges.scala 447:17 452:15]
  assign auto_mem_out_a_bits_mask = {x1_a_bits_a_mask_hi,x1_a_bits_a_mask_lo}; // @[Cat.scala 33:92]
  assign auto_mem_out_d_ready = loader_io_cache_block_in_ready; // @[Nodes.scala 1212:84 CScratchpad.scala 180:19]
  assign loader_clock = clock;
  assign loader_reset = reset;
  assign loader_io_cache_block_in_valid = auto_mem_out_d_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign loader_io_cache_block_in_bits_len = _GEN_235[6:0];
  always @(posedge clock) begin
    if (reset) begin // @[CScratchpad.scala 102:37]
      mem_tx_state <= 2'h0; // @[CScratchpad.scala 102:37]
    end else if (!(2'h0 == mem_tx_state)) begin // @[CScratchpad.scala 138:24]
      if (2'h1 == mem_tx_state) begin // @[CScratchpad.scala 138:24]
        if (_T_13) begin // @[CScratchpad.scala 152:28]
          mem_tx_state <= _GEN_56;
        end
      end else if (2'h2 == mem_tx_state) begin // @[CScratchpad.scala 138:24]
        mem_tx_state <= _GEN_109;
      end
    end
    reqIdleBits_0 <= reset | _GEN_494; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_1 <= reset | _GEN_495; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_2 <= reset | _GEN_496; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_3 <= reset | _GEN_497; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_4 <= reset | _GEN_498; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_5 <= reset | _GEN_499; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_6 <= reset | _GEN_500; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_7 <= reset | _GEN_501; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_8 <= reset | _GEN_502; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_9 <= reset | _GEN_503; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_10 <= reset | _GEN_504; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_11 <= reset | _GEN_505; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_12 <= reset | _GEN_506; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_13 <= reset | _GEN_507; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_14 <= reset | _GEN_508; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_15 <= reset | _GEN_509; // @[CScratchpad.scala 110:{36,36}]
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h0 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_0_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_0_memoryLength <= _GEN_203;
      end
    end else begin
      req_cache_0_memoryLength <= _GEN_203;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h1 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_1_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_1_memoryLength <= _GEN_204;
      end
    end else begin
      req_cache_1_memoryLength <= _GEN_204;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h2 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_2_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_2_memoryLength <= _GEN_205;
      end
    end else begin
      req_cache_2_memoryLength <= _GEN_205;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h3 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_3_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_3_memoryLength <= _GEN_206;
      end
    end else begin
      req_cache_3_memoryLength <= _GEN_206;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h4 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_4_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_4_memoryLength <= _GEN_207;
      end
    end else begin
      req_cache_4_memoryLength <= _GEN_207;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h5 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_5_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_5_memoryLength <= _GEN_208;
      end
    end else begin
      req_cache_5_memoryLength <= _GEN_208;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h6 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_6_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_6_memoryLength <= _GEN_209;
      end
    end else begin
      req_cache_6_memoryLength <= _GEN_209;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h7 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_7_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_7_memoryLength <= _GEN_210;
      end
    end else begin
      req_cache_7_memoryLength <= _GEN_210;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h8 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_8_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_8_memoryLength <= _GEN_211;
      end
    end else begin
      req_cache_8_memoryLength <= _GEN_211;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h9 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_9_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_9_memoryLength <= _GEN_212;
      end
    end else begin
      req_cache_9_memoryLength <= _GEN_212;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'ha == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_10_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_10_memoryLength <= _GEN_213;
      end
    end else begin
      req_cache_10_memoryLength <= _GEN_213;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'hb == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_11_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_11_memoryLength <= _GEN_214;
      end
    end else begin
      req_cache_11_memoryLength <= _GEN_214;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'hc == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_12_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_12_memoryLength <= _GEN_215;
      end
    end else begin
      req_cache_12_memoryLength <= _GEN_215;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'hd == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_13_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_13_memoryLength <= _GEN_216;
      end
    end else begin
      req_cache_13_memoryLength <= _GEN_216;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'he == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_14_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_14_memoryLength <= _GEN_217;
      end
    end else begin
      req_cache_14_memoryLength <= _GEN_217;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'hf == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_15_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_15_memoryLength <= _GEN_218;
      end
    end else begin
      req_cache_15_memoryLength <= _GEN_218;
    end
    if (!(2'h0 == mem_tx_state)) begin // @[CScratchpad.scala 138:24]
      if (2'h1 == mem_tx_state) begin // @[CScratchpad.scala 138:24]
        if (_T_13) begin // @[CScratchpad.scala 152:28]
          totalTx_memoryAddress <= _totalTx_memoryAddress_T_1; // @[CScratchpad.scala 158:31]
        end
      end
    end
    if (!(2'h0 == mem_tx_state)) begin // @[CScratchpad.scala 138:24]
      if (2'h1 == mem_tx_state) begin // @[CScratchpad.scala 138:24]
        if (_T_13) begin // @[CScratchpad.scala 152:28]
          totalTx_memoryLength <= _totalTx_memoryLength_T_1; // @[CScratchpad.scala 156:30]
        end
      end
    end
  end
endmodule
module CScratchpadPackedSubwordLoader_2(
  input        clock,
  input        reset,
  output       io_cache_block_in_ready,
  input        io_cache_block_in_valid,
  input  [6:0] io_cache_block_in_bits_len,
  output       io_sp_write_out_valid
);
  reg [6:0] lenRemainingFromReq; // @[CScratchpadPackedSubwordLoader.scala 18:32]
  reg  state; // @[CScratchpadPackedSubwordLoader.scala 21:22]
  wire  _io_cache_block_in_ready_T = ~state; // @[CScratchpadPackedSubwordLoader.scala 22:36]
  wire  _T_1 = io_cache_block_in_ready & io_cache_block_in_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_0 = _T_1 | state; // @[CScratchpadPackedSubwordLoader.scala 34:36 35:15 21:22]
  wire [6:0] _lenRemainingFromReq_T_1 = lenRemainingFromReq - 7'h20; // @[CScratchpadPackedSubwordLoader.scala 53:54]
  wire  _GEN_6 = lenRemainingFromReq == 7'h20 ? 1'h0 : state; // @[CScratchpadPackedSubwordLoader.scala 54:60 55:19 21:22]
  assign io_cache_block_in_ready = ~state; // @[CScratchpadPackedSubwordLoader.scala 22:36]
  assign io_sp_write_out_valid = _io_cache_block_in_ready_T ? 1'h0 : state; // @[CScratchpadPackedSubwordLoader.scala 32:17 24:25]
  always @(posedge clock) begin
    if (_io_cache_block_in_ready_T) begin // @[CScratchpadPackedSubwordLoader.scala 32:17]
      if (_T_1) begin // @[CScratchpadPackedSubwordLoader.scala 34:36]
        lenRemainingFromReq <= io_cache_block_in_bits_len; // @[CScratchpadPackedSubwordLoader.scala 38:29]
      end
    end else if (state) begin // @[CScratchpadPackedSubwordLoader.scala 32:17]
      if (io_sp_write_out_valid) begin // @[CScratchpadPackedSubwordLoader.scala 48:34]
        lenRemainingFromReq <= _lenRemainingFromReq_T_1;
      end
    end
    if (reset) begin // @[CScratchpadPackedSubwordLoader.scala 21:22]
      state <= 1'h0; // @[CScratchpadPackedSubwordLoader.scala 21:22]
    end else if (_io_cache_block_in_ready_T) begin // @[CScratchpadPackedSubwordLoader.scala 32:17]
      state <= _GEN_0;
    end else if (state) begin // @[CScratchpadPackedSubwordLoader.scala 32:17]
      if (io_sp_write_out_valid) begin // @[CScratchpadPackedSubwordLoader.scala 48:34]
        state <= _GEN_6;
      end
    end
  end
endmodule
module CScratchpad_2(
  input         clock,
  input         reset,
  input         auto_mem_out_a_ready,
  output        auto_mem_out_a_valid,
  output [2:0]  auto_mem_out_a_bits_size,
  output [3:0]  auto_mem_out_a_bits_source,
  output [33:0] auto_mem_out_a_bits_address,
  output [63:0] auto_mem_out_a_bits_mask,
  output        auto_mem_out_d_ready,
  input         auto_mem_out_d_valid,
  input  [3:0]  auto_mem_out_d_bits_source
);
  wire  loader_clock; // @[CScratchpad.scala 94:30]
  wire  loader_reset; // @[CScratchpad.scala 94:30]
  wire  loader_io_cache_block_in_ready; // @[CScratchpad.scala 94:30]
  wire  loader_io_cache_block_in_valid; // @[CScratchpad.scala 94:30]
  wire [6:0] loader_io_cache_block_in_bits_len; // @[CScratchpad.scala 94:30]
  wire  loader_io_sp_write_out_valid; // @[CScratchpad.scala 94:30]
  reg [1:0] mem_tx_state; // @[CScratchpad.scala 102:37]
  reg  reqIdleBits_0; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_1; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_2; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_3; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_4; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_5; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_6; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_7; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_8; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_9; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_10; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_11; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_12; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_13; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_14; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_15; // @[CScratchpad.scala 110:36]
  wire  reqAvailable = reqIdleBits_0 | reqIdleBits_1 | reqIdleBits_2 | reqIdleBits_3 | reqIdleBits_4 | reqIdleBits_5 |
    reqIdleBits_6 | reqIdleBits_7 | reqIdleBits_8 | reqIdleBits_9 | reqIdleBits_10 | reqIdleBits_11 | reqIdleBits_12 |
    reqIdleBits_13 | reqIdleBits_14 | reqIdleBits_15; // @[CScratchpad.scala 111:51]
  wire [3:0] _reqChosen_T = reqIdleBits_14 ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_1 = reqIdleBits_13 ? 4'hd : _reqChosen_T; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_2 = reqIdleBits_12 ? 4'hc : _reqChosen_T_1; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_3 = reqIdleBits_11 ? 4'hb : _reqChosen_T_2; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_4 = reqIdleBits_10 ? 4'ha : _reqChosen_T_3; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_5 = reqIdleBits_9 ? 4'h9 : _reqChosen_T_4; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_6 = reqIdleBits_8 ? 4'h8 : _reqChosen_T_5; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_7 = reqIdleBits_7 ? 4'h7 : _reqChosen_T_6; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_8 = reqIdleBits_6 ? 4'h6 : _reqChosen_T_7; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_9 = reqIdleBits_5 ? 4'h5 : _reqChosen_T_8; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_10 = reqIdleBits_4 ? 4'h4 : _reqChosen_T_9; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_11 = reqIdleBits_3 ? 4'h3 : _reqChosen_T_10; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_12 = reqIdleBits_2 ? 4'h2 : _reqChosen_T_11; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_13 = reqIdleBits_1 ? 4'h1 : _reqChosen_T_12; // @[Mux.scala 47:70]
  wire [3:0] reqChosen = reqIdleBits_0 ? 4'h0 : _reqChosen_T_13; // @[Mux.scala 47:70]
  reg [15:0] req_cache_0_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_1_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_2_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_3_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_4_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_5_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_6_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_7_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_8_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_9_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_10_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_11_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_12_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_13_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_14_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_15_memoryLength; // @[CScratchpad.scala 114:30]
  reg [33:0] totalTx_memoryAddress; // @[CScratchpad.scala 124:28]
  reg [33:0] totalTx_memoryLength; // @[CScratchpad.scala 124:28]
  wire  isBelowLimit = totalTx_memoryLength <= 34'h40; // @[CScratchpad.scala 149:47]
  wire [1:0] txEmitLengthLg_hi = totalTx_memoryLength[33:32]; // @[OneHot.scala 30:18]
  wire  _txEmitLengthLg_T = |txEmitLengthLg_hi; // @[OneHot.scala 32:14]
  wire [31:0] txEmitLengthLg_lo = totalTx_memoryLength[31:0]; // @[OneHot.scala 31:18]
  wire [31:0] _GEN_569 = {{30'd0}, txEmitLengthLg_hi}; // @[OneHot.scala 32:28]
  wire [31:0] _txEmitLengthLg_T_1 = _GEN_569 | txEmitLengthLg_lo; // @[OneHot.scala 32:28]
  wire [15:0] txEmitLengthLg_hi_1 = _txEmitLengthLg_T_1[31:16]; // @[OneHot.scala 30:18]
  wire  _txEmitLengthLg_T_2 = |txEmitLengthLg_hi_1; // @[OneHot.scala 32:14]
  wire [15:0] txEmitLengthLg_lo_1 = _txEmitLengthLg_T_1[15:0]; // @[OneHot.scala 31:18]
  wire [15:0] _txEmitLengthLg_T_3 = txEmitLengthLg_hi_1 | txEmitLengthLg_lo_1; // @[OneHot.scala 32:28]
  wire [7:0] txEmitLengthLg_hi_2 = _txEmitLengthLg_T_3[15:8]; // @[OneHot.scala 30:18]
  wire  _txEmitLengthLg_T_4 = |txEmitLengthLg_hi_2; // @[OneHot.scala 32:14]
  wire [7:0] txEmitLengthLg_lo_2 = _txEmitLengthLg_T_3[7:0]; // @[OneHot.scala 31:18]
  wire [7:0] _txEmitLengthLg_T_5 = txEmitLengthLg_hi_2 | txEmitLengthLg_lo_2; // @[OneHot.scala 32:28]
  wire [3:0] txEmitLengthLg_hi_3 = _txEmitLengthLg_T_5[7:4]; // @[OneHot.scala 30:18]
  wire  _txEmitLengthLg_T_6 = |txEmitLengthLg_hi_3; // @[OneHot.scala 32:14]
  wire [3:0] txEmitLengthLg_lo_3 = _txEmitLengthLg_T_5[3:0]; // @[OneHot.scala 31:18]
  wire [3:0] _txEmitLengthLg_T_7 = txEmitLengthLg_hi_3 | txEmitLengthLg_lo_3; // @[OneHot.scala 32:28]
  wire [1:0] txEmitLengthLg_hi_4 = _txEmitLengthLg_T_7[3:2]; // @[OneHot.scala 30:18]
  wire  _txEmitLengthLg_T_8 = |txEmitLengthLg_hi_4; // @[OneHot.scala 32:14]
  wire [1:0] txEmitLengthLg_lo_4 = _txEmitLengthLg_T_7[1:0]; // @[OneHot.scala 31:18]
  wire [1:0] _txEmitLengthLg_T_9 = txEmitLengthLg_hi_4 | txEmitLengthLg_lo_4; // @[OneHot.scala 32:28]
  wire [5:0] _txEmitLengthLg_T_15 = {_txEmitLengthLg_T,_txEmitLengthLg_T_2,_txEmitLengthLg_T_4,_txEmitLengthLg_T_6,
    _txEmitLengthLg_T_8,_txEmitLengthLg_T_9[1]}; // @[Cat.scala 33:92]
  wire [5:0] _txEmitLengthLg_T_16 = isBelowLimit ? _txEmitLengthLg_T_15 : 6'h6; // @[CScratchpad.scala 150:28]
  wire [5:0] _GEN_111 = 2'h1 == mem_tx_state ? _txEmitLengthLg_T_16 : 6'h0; // @[CScratchpad.scala 131:18 138:24 150:22]
  wire [5:0] _GEN_169 = 2'h0 == mem_tx_state ? 6'h0 : _GEN_111; // @[CScratchpad.scala 131:18 138:24]
  wire [3:0] txEmitLengthLg = _GEN_169[3:0]; // @[CScratchpad.scala 130:36]
  wire [5:0] _x1_a_bits_a_mask_sizeOH_T = {{2'd0}, txEmitLengthLg}; // @[Misc.scala 201:34]
  wire [2:0] x1_a_bits_a_mask_sizeOH_shiftAmount = _x1_a_bits_a_mask_sizeOH_T[2:0]; // @[OneHot.scala 63:49]
  wire [7:0] _x1_a_bits_a_mask_sizeOH_T_1 = 8'h1 << x1_a_bits_a_mask_sizeOH_shiftAmount; // @[OneHot.scala 64:12]
  wire [5:0] x1_a_bits_a_mask_sizeOH = _x1_a_bits_a_mask_sizeOH_T_1[5:0] | 6'h1; // @[Misc.scala 201:81]
  wire  _x1_a_bits_a_mask_T = txEmitLengthLg >= 4'h6; // @[Misc.scala 205:21]
  wire  x1_a_bits_a_mask_size = x1_a_bits_a_mask_sizeOH[5]; // @[Misc.scala 208:26]
  wire  x1_a_bits_a_mask_bit = totalTx_memoryAddress[5]; // @[Misc.scala 209:26]
  wire  x1_a_bits_a_mask_nbit = ~x1_a_bits_a_mask_bit; // @[Misc.scala 210:20]
  wire  x1_a_bits_a_mask_acc = _x1_a_bits_a_mask_T | x1_a_bits_a_mask_size & x1_a_bits_a_mask_nbit; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_acc_1 = _x1_a_bits_a_mask_T | x1_a_bits_a_mask_size & x1_a_bits_a_mask_bit; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_size_1 = x1_a_bits_a_mask_sizeOH[4]; // @[Misc.scala 208:26]
  wire  x1_a_bits_a_mask_bit_1 = totalTx_memoryAddress[4]; // @[Misc.scala 209:26]
  wire  x1_a_bits_a_mask_nbit_1 = ~x1_a_bits_a_mask_bit_1; // @[Misc.scala 210:20]
  wire  x1_a_bits_a_mask_eq_2 = x1_a_bits_a_mask_nbit & x1_a_bits_a_mask_nbit_1; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_2 = x1_a_bits_a_mask_acc | x1_a_bits_a_mask_size_1 & x1_a_bits_a_mask_eq_2; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_3 = x1_a_bits_a_mask_nbit & x1_a_bits_a_mask_bit_1; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_3 = x1_a_bits_a_mask_acc | x1_a_bits_a_mask_size_1 & x1_a_bits_a_mask_eq_3; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_4 = x1_a_bits_a_mask_bit & x1_a_bits_a_mask_nbit_1; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_4 = x1_a_bits_a_mask_acc_1 | x1_a_bits_a_mask_size_1 & x1_a_bits_a_mask_eq_4; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_5 = x1_a_bits_a_mask_bit & x1_a_bits_a_mask_bit_1; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_5 = x1_a_bits_a_mask_acc_1 | x1_a_bits_a_mask_size_1 & x1_a_bits_a_mask_eq_5; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_size_2 = x1_a_bits_a_mask_sizeOH[3]; // @[Misc.scala 208:26]
  wire  x1_a_bits_a_mask_bit_2 = totalTx_memoryAddress[3]; // @[Misc.scala 209:26]
  wire  x1_a_bits_a_mask_nbit_2 = ~x1_a_bits_a_mask_bit_2; // @[Misc.scala 210:20]
  wire  x1_a_bits_a_mask_eq_6 = x1_a_bits_a_mask_eq_2 & x1_a_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_6 = x1_a_bits_a_mask_acc_2 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_6; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_7 = x1_a_bits_a_mask_eq_2 & x1_a_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_7 = x1_a_bits_a_mask_acc_2 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_7; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_8 = x1_a_bits_a_mask_eq_3 & x1_a_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_8 = x1_a_bits_a_mask_acc_3 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_8; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_9 = x1_a_bits_a_mask_eq_3 & x1_a_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_9 = x1_a_bits_a_mask_acc_3 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_9; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_10 = x1_a_bits_a_mask_eq_4 & x1_a_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_10 = x1_a_bits_a_mask_acc_4 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_10; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_11 = x1_a_bits_a_mask_eq_4 & x1_a_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_11 = x1_a_bits_a_mask_acc_4 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_11; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_12 = x1_a_bits_a_mask_eq_5 & x1_a_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_12 = x1_a_bits_a_mask_acc_5 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_12; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_13 = x1_a_bits_a_mask_eq_5 & x1_a_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_13 = x1_a_bits_a_mask_acc_5 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_13; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_size_3 = x1_a_bits_a_mask_sizeOH[2]; // @[Misc.scala 208:26]
  wire  x1_a_bits_a_mask_bit_3 = totalTx_memoryAddress[2]; // @[Misc.scala 209:26]
  wire  x1_a_bits_a_mask_nbit_3 = ~x1_a_bits_a_mask_bit_3; // @[Misc.scala 210:20]
  wire  x1_a_bits_a_mask_eq_14 = x1_a_bits_a_mask_eq_6 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_14 = x1_a_bits_a_mask_acc_6 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_14; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_15 = x1_a_bits_a_mask_eq_6 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_15 = x1_a_bits_a_mask_acc_6 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_15; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_16 = x1_a_bits_a_mask_eq_7 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_16 = x1_a_bits_a_mask_acc_7 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_16; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_17 = x1_a_bits_a_mask_eq_7 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_17 = x1_a_bits_a_mask_acc_7 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_17; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_18 = x1_a_bits_a_mask_eq_8 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_18 = x1_a_bits_a_mask_acc_8 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_18; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_19 = x1_a_bits_a_mask_eq_8 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_19 = x1_a_bits_a_mask_acc_8 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_19; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_20 = x1_a_bits_a_mask_eq_9 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_20 = x1_a_bits_a_mask_acc_9 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_20; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_21 = x1_a_bits_a_mask_eq_9 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_21 = x1_a_bits_a_mask_acc_9 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_21; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_22 = x1_a_bits_a_mask_eq_10 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_22 = x1_a_bits_a_mask_acc_10 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_22; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_23 = x1_a_bits_a_mask_eq_10 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_23 = x1_a_bits_a_mask_acc_10 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_23; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_24 = x1_a_bits_a_mask_eq_11 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_24 = x1_a_bits_a_mask_acc_11 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_24; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_25 = x1_a_bits_a_mask_eq_11 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_25 = x1_a_bits_a_mask_acc_11 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_25; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_26 = x1_a_bits_a_mask_eq_12 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_26 = x1_a_bits_a_mask_acc_12 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_26; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_27 = x1_a_bits_a_mask_eq_12 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_27 = x1_a_bits_a_mask_acc_12 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_27; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_28 = x1_a_bits_a_mask_eq_13 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_28 = x1_a_bits_a_mask_acc_13 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_28; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_29 = x1_a_bits_a_mask_eq_13 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_29 = x1_a_bits_a_mask_acc_13 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_29; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_size_4 = x1_a_bits_a_mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  x1_a_bits_a_mask_bit_4 = totalTx_memoryAddress[1]; // @[Misc.scala 209:26]
  wire  x1_a_bits_a_mask_nbit_4 = ~x1_a_bits_a_mask_bit_4; // @[Misc.scala 210:20]
  wire  x1_a_bits_a_mask_eq_30 = x1_a_bits_a_mask_eq_14 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_30 = x1_a_bits_a_mask_acc_14 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_30; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_31 = x1_a_bits_a_mask_eq_14 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_31 = x1_a_bits_a_mask_acc_14 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_31; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_32 = x1_a_bits_a_mask_eq_15 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_32 = x1_a_bits_a_mask_acc_15 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_32; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_33 = x1_a_bits_a_mask_eq_15 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_33 = x1_a_bits_a_mask_acc_15 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_33; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_34 = x1_a_bits_a_mask_eq_16 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_34 = x1_a_bits_a_mask_acc_16 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_34; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_35 = x1_a_bits_a_mask_eq_16 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_35 = x1_a_bits_a_mask_acc_16 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_35; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_36 = x1_a_bits_a_mask_eq_17 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_36 = x1_a_bits_a_mask_acc_17 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_36; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_37 = x1_a_bits_a_mask_eq_17 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_37 = x1_a_bits_a_mask_acc_17 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_37; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_38 = x1_a_bits_a_mask_eq_18 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_38 = x1_a_bits_a_mask_acc_18 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_38; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_39 = x1_a_bits_a_mask_eq_18 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_39 = x1_a_bits_a_mask_acc_18 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_39; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_40 = x1_a_bits_a_mask_eq_19 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_40 = x1_a_bits_a_mask_acc_19 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_40; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_41 = x1_a_bits_a_mask_eq_19 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_41 = x1_a_bits_a_mask_acc_19 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_41; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_42 = x1_a_bits_a_mask_eq_20 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_42 = x1_a_bits_a_mask_acc_20 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_42; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_43 = x1_a_bits_a_mask_eq_20 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_43 = x1_a_bits_a_mask_acc_20 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_43; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_44 = x1_a_bits_a_mask_eq_21 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_44 = x1_a_bits_a_mask_acc_21 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_44; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_45 = x1_a_bits_a_mask_eq_21 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_45 = x1_a_bits_a_mask_acc_21 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_45; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_46 = x1_a_bits_a_mask_eq_22 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_46 = x1_a_bits_a_mask_acc_22 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_46; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_47 = x1_a_bits_a_mask_eq_22 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_47 = x1_a_bits_a_mask_acc_22 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_47; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_48 = x1_a_bits_a_mask_eq_23 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_48 = x1_a_bits_a_mask_acc_23 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_48; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_49 = x1_a_bits_a_mask_eq_23 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_49 = x1_a_bits_a_mask_acc_23 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_49; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_50 = x1_a_bits_a_mask_eq_24 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_50 = x1_a_bits_a_mask_acc_24 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_50; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_51 = x1_a_bits_a_mask_eq_24 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_51 = x1_a_bits_a_mask_acc_24 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_51; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_52 = x1_a_bits_a_mask_eq_25 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_52 = x1_a_bits_a_mask_acc_25 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_52; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_53 = x1_a_bits_a_mask_eq_25 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_53 = x1_a_bits_a_mask_acc_25 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_53; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_54 = x1_a_bits_a_mask_eq_26 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_54 = x1_a_bits_a_mask_acc_26 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_54; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_55 = x1_a_bits_a_mask_eq_26 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_55 = x1_a_bits_a_mask_acc_26 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_55; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_56 = x1_a_bits_a_mask_eq_27 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_56 = x1_a_bits_a_mask_acc_27 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_56; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_57 = x1_a_bits_a_mask_eq_27 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_57 = x1_a_bits_a_mask_acc_27 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_57; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_58 = x1_a_bits_a_mask_eq_28 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_58 = x1_a_bits_a_mask_acc_28 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_58; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_59 = x1_a_bits_a_mask_eq_28 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_59 = x1_a_bits_a_mask_acc_28 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_59; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_60 = x1_a_bits_a_mask_eq_29 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_60 = x1_a_bits_a_mask_acc_29 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_60; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_61 = x1_a_bits_a_mask_eq_29 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_61 = x1_a_bits_a_mask_acc_29 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_61; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_size_5 = x1_a_bits_a_mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  x1_a_bits_a_mask_bit_5 = totalTx_memoryAddress[0]; // @[Misc.scala 209:26]
  wire  x1_a_bits_a_mask_nbit_5 = ~x1_a_bits_a_mask_bit_5; // @[Misc.scala 210:20]
  wire  x1_a_bits_a_mask_eq_62 = x1_a_bits_a_mask_eq_30 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_62 = x1_a_bits_a_mask_acc_30 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_62; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_63 = x1_a_bits_a_mask_eq_30 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_63 = x1_a_bits_a_mask_acc_30 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_63; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_64 = x1_a_bits_a_mask_eq_31 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_64 = x1_a_bits_a_mask_acc_31 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_64; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_65 = x1_a_bits_a_mask_eq_31 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_65 = x1_a_bits_a_mask_acc_31 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_65; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_66 = x1_a_bits_a_mask_eq_32 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_66 = x1_a_bits_a_mask_acc_32 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_66; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_67 = x1_a_bits_a_mask_eq_32 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_67 = x1_a_bits_a_mask_acc_32 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_67; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_68 = x1_a_bits_a_mask_eq_33 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_68 = x1_a_bits_a_mask_acc_33 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_68; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_69 = x1_a_bits_a_mask_eq_33 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_69 = x1_a_bits_a_mask_acc_33 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_69; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_70 = x1_a_bits_a_mask_eq_34 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_70 = x1_a_bits_a_mask_acc_34 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_70; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_71 = x1_a_bits_a_mask_eq_34 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_71 = x1_a_bits_a_mask_acc_34 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_71; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_72 = x1_a_bits_a_mask_eq_35 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_72 = x1_a_bits_a_mask_acc_35 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_72; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_73 = x1_a_bits_a_mask_eq_35 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_73 = x1_a_bits_a_mask_acc_35 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_73; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_74 = x1_a_bits_a_mask_eq_36 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_74 = x1_a_bits_a_mask_acc_36 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_74; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_75 = x1_a_bits_a_mask_eq_36 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_75 = x1_a_bits_a_mask_acc_36 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_75; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_76 = x1_a_bits_a_mask_eq_37 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_76 = x1_a_bits_a_mask_acc_37 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_76; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_77 = x1_a_bits_a_mask_eq_37 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_77 = x1_a_bits_a_mask_acc_37 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_77; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_78 = x1_a_bits_a_mask_eq_38 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_78 = x1_a_bits_a_mask_acc_38 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_78; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_79 = x1_a_bits_a_mask_eq_38 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_79 = x1_a_bits_a_mask_acc_38 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_79; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_80 = x1_a_bits_a_mask_eq_39 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_80 = x1_a_bits_a_mask_acc_39 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_80; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_81 = x1_a_bits_a_mask_eq_39 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_81 = x1_a_bits_a_mask_acc_39 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_81; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_82 = x1_a_bits_a_mask_eq_40 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_82 = x1_a_bits_a_mask_acc_40 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_82; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_83 = x1_a_bits_a_mask_eq_40 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_83 = x1_a_bits_a_mask_acc_40 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_83; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_84 = x1_a_bits_a_mask_eq_41 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_84 = x1_a_bits_a_mask_acc_41 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_84; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_85 = x1_a_bits_a_mask_eq_41 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_85 = x1_a_bits_a_mask_acc_41 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_85; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_86 = x1_a_bits_a_mask_eq_42 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_86 = x1_a_bits_a_mask_acc_42 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_86; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_87 = x1_a_bits_a_mask_eq_42 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_87 = x1_a_bits_a_mask_acc_42 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_87; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_88 = x1_a_bits_a_mask_eq_43 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_88 = x1_a_bits_a_mask_acc_43 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_88; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_89 = x1_a_bits_a_mask_eq_43 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_89 = x1_a_bits_a_mask_acc_43 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_89; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_90 = x1_a_bits_a_mask_eq_44 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_90 = x1_a_bits_a_mask_acc_44 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_90; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_91 = x1_a_bits_a_mask_eq_44 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_91 = x1_a_bits_a_mask_acc_44 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_91; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_92 = x1_a_bits_a_mask_eq_45 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_92 = x1_a_bits_a_mask_acc_45 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_92; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_93 = x1_a_bits_a_mask_eq_45 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_93 = x1_a_bits_a_mask_acc_45 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_93; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_94 = x1_a_bits_a_mask_eq_46 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_94 = x1_a_bits_a_mask_acc_46 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_94; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_95 = x1_a_bits_a_mask_eq_46 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_95 = x1_a_bits_a_mask_acc_46 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_95; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_96 = x1_a_bits_a_mask_eq_47 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_96 = x1_a_bits_a_mask_acc_47 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_96; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_97 = x1_a_bits_a_mask_eq_47 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_97 = x1_a_bits_a_mask_acc_47 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_97; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_98 = x1_a_bits_a_mask_eq_48 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_98 = x1_a_bits_a_mask_acc_48 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_98; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_99 = x1_a_bits_a_mask_eq_48 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_99 = x1_a_bits_a_mask_acc_48 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_99; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_100 = x1_a_bits_a_mask_eq_49 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_100 = x1_a_bits_a_mask_acc_49 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_100; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_101 = x1_a_bits_a_mask_eq_49 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_101 = x1_a_bits_a_mask_acc_49 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_101; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_102 = x1_a_bits_a_mask_eq_50 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_102 = x1_a_bits_a_mask_acc_50 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_102; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_103 = x1_a_bits_a_mask_eq_50 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_103 = x1_a_bits_a_mask_acc_50 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_103; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_104 = x1_a_bits_a_mask_eq_51 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_104 = x1_a_bits_a_mask_acc_51 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_104; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_105 = x1_a_bits_a_mask_eq_51 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_105 = x1_a_bits_a_mask_acc_51 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_105; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_106 = x1_a_bits_a_mask_eq_52 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_106 = x1_a_bits_a_mask_acc_52 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_106; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_107 = x1_a_bits_a_mask_eq_52 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_107 = x1_a_bits_a_mask_acc_52 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_107; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_108 = x1_a_bits_a_mask_eq_53 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_108 = x1_a_bits_a_mask_acc_53 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_108; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_109 = x1_a_bits_a_mask_eq_53 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_109 = x1_a_bits_a_mask_acc_53 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_109; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_110 = x1_a_bits_a_mask_eq_54 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_110 = x1_a_bits_a_mask_acc_54 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_110; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_111 = x1_a_bits_a_mask_eq_54 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_111 = x1_a_bits_a_mask_acc_54 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_111; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_112 = x1_a_bits_a_mask_eq_55 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_112 = x1_a_bits_a_mask_acc_55 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_112; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_113 = x1_a_bits_a_mask_eq_55 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_113 = x1_a_bits_a_mask_acc_55 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_113; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_114 = x1_a_bits_a_mask_eq_56 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_114 = x1_a_bits_a_mask_acc_56 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_114; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_115 = x1_a_bits_a_mask_eq_56 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_115 = x1_a_bits_a_mask_acc_56 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_115; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_116 = x1_a_bits_a_mask_eq_57 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_116 = x1_a_bits_a_mask_acc_57 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_116; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_117 = x1_a_bits_a_mask_eq_57 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_117 = x1_a_bits_a_mask_acc_57 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_117; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_118 = x1_a_bits_a_mask_eq_58 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_118 = x1_a_bits_a_mask_acc_58 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_118; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_119 = x1_a_bits_a_mask_eq_58 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_119 = x1_a_bits_a_mask_acc_58 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_119; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_120 = x1_a_bits_a_mask_eq_59 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_120 = x1_a_bits_a_mask_acc_59 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_120; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_121 = x1_a_bits_a_mask_eq_59 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_121 = x1_a_bits_a_mask_acc_59 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_121; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_122 = x1_a_bits_a_mask_eq_60 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_122 = x1_a_bits_a_mask_acc_60 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_122; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_123 = x1_a_bits_a_mask_eq_60 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_123 = x1_a_bits_a_mask_acc_60 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_123; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_124 = x1_a_bits_a_mask_eq_61 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_124 = x1_a_bits_a_mask_acc_61 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_124; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_125 = x1_a_bits_a_mask_eq_61 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_125 = x1_a_bits_a_mask_acc_61 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_125; // @[Misc.scala 214:29]
  wire [7:0] x1_a_bits_a_mask_lo_lo_lo = {x1_a_bits_a_mask_acc_69,x1_a_bits_a_mask_acc_68,x1_a_bits_a_mask_acc_67,
    x1_a_bits_a_mask_acc_66,x1_a_bits_a_mask_acc_65,x1_a_bits_a_mask_acc_64,x1_a_bits_a_mask_acc_63,
    x1_a_bits_a_mask_acc_62}; // @[Cat.scala 33:92]
  wire [15:0] x1_a_bits_a_mask_lo_lo = {x1_a_bits_a_mask_acc_77,x1_a_bits_a_mask_acc_76,x1_a_bits_a_mask_acc_75,
    x1_a_bits_a_mask_acc_74,x1_a_bits_a_mask_acc_73,x1_a_bits_a_mask_acc_72,x1_a_bits_a_mask_acc_71,
    x1_a_bits_a_mask_acc_70,x1_a_bits_a_mask_lo_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] x1_a_bits_a_mask_lo_hi_lo = {x1_a_bits_a_mask_acc_85,x1_a_bits_a_mask_acc_84,x1_a_bits_a_mask_acc_83,
    x1_a_bits_a_mask_acc_82,x1_a_bits_a_mask_acc_81,x1_a_bits_a_mask_acc_80,x1_a_bits_a_mask_acc_79,
    x1_a_bits_a_mask_acc_78}; // @[Cat.scala 33:92]
  wire [31:0] x1_a_bits_a_mask_lo = {x1_a_bits_a_mask_acc_93,x1_a_bits_a_mask_acc_92,x1_a_bits_a_mask_acc_91,
    x1_a_bits_a_mask_acc_90,x1_a_bits_a_mask_acc_89,x1_a_bits_a_mask_acc_88,x1_a_bits_a_mask_acc_87,
    x1_a_bits_a_mask_acc_86,x1_a_bits_a_mask_lo_hi_lo,x1_a_bits_a_mask_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] x1_a_bits_a_mask_hi_lo_lo = {x1_a_bits_a_mask_acc_101,x1_a_bits_a_mask_acc_100,x1_a_bits_a_mask_acc_99,
    x1_a_bits_a_mask_acc_98,x1_a_bits_a_mask_acc_97,x1_a_bits_a_mask_acc_96,x1_a_bits_a_mask_acc_95,
    x1_a_bits_a_mask_acc_94}; // @[Cat.scala 33:92]
  wire [15:0] x1_a_bits_a_mask_hi_lo = {x1_a_bits_a_mask_acc_109,x1_a_bits_a_mask_acc_108,x1_a_bits_a_mask_acc_107,
    x1_a_bits_a_mask_acc_106,x1_a_bits_a_mask_acc_105,x1_a_bits_a_mask_acc_104,x1_a_bits_a_mask_acc_103,
    x1_a_bits_a_mask_acc_102,x1_a_bits_a_mask_hi_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] x1_a_bits_a_mask_hi_hi_lo = {x1_a_bits_a_mask_acc_117,x1_a_bits_a_mask_acc_116,x1_a_bits_a_mask_acc_115,
    x1_a_bits_a_mask_acc_114,x1_a_bits_a_mask_acc_113,x1_a_bits_a_mask_acc_112,x1_a_bits_a_mask_acc_111,
    x1_a_bits_a_mask_acc_110}; // @[Cat.scala 33:92]
  wire [31:0] x1_a_bits_a_mask_hi = {x1_a_bits_a_mask_acc_125,x1_a_bits_a_mask_acc_124,x1_a_bits_a_mask_acc_123,
    x1_a_bits_a_mask_acc_122,x1_a_bits_a_mask_acc_121,x1_a_bits_a_mask_acc_120,x1_a_bits_a_mask_acc_119,
    x1_a_bits_a_mask_acc_118,x1_a_bits_a_mask_hi_hi_lo,x1_a_bits_a_mask_hi_lo}; // @[Cat.scala 33:92]
  wire  _GEN_112 = 2'h1 == mem_tx_state ? reqAvailable : mem_tx_state == 2'h1; // @[CScratchpad.scala 136:19 138:24 151:23]
  wire  mem_out_a_valid = 2'h0 == mem_tx_state ? mem_tx_state == 2'h1 : _GEN_112; // @[CScratchpad.scala 136:19 138:24]
  wire  _T_13 = auto_mem_out_a_ready & mem_out_a_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_8 = 4'h0 == reqChosen ? 1'h0 : reqIdleBits_0; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_9 = 4'h1 == reqChosen ? 1'h0 : reqIdleBits_1; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_10 = 4'h2 == reqChosen ? 1'h0 : reqIdleBits_2; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_11 = 4'h3 == reqChosen ? 1'h0 : reqIdleBits_3; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_12 = 4'h4 == reqChosen ? 1'h0 : reqIdleBits_4; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_13 = 4'h5 == reqChosen ? 1'h0 : reqIdleBits_5; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_14 = 4'h6 == reqChosen ? 1'h0 : reqIdleBits_6; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_15 = 4'h7 == reqChosen ? 1'h0 : reqIdleBits_7; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_16 = 4'h8 == reqChosen ? 1'h0 : reqIdleBits_8; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_17 = 4'h9 == reqChosen ? 1'h0 : reqIdleBits_9; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_18 = 4'ha == reqChosen ? 1'h0 : reqIdleBits_10; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_19 = 4'hb == reqChosen ? 1'h0 : reqIdleBits_11; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_20 = 4'hc == reqChosen ? 1'h0 : reqIdleBits_12; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_21 = 4'hd == reqChosen ? 1'h0 : reqIdleBits_13; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_22 = 4'he == reqChosen ? 1'h0 : reqIdleBits_14; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_23 = 4'hf == reqChosen ? 1'h0 : reqIdleBits_15; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire [33:0] _req_cache_memoryLength_T = isBelowLimit ? totalTx_memoryLength : 34'h40; // @[CScratchpad.scala 155:49]
  wire [15:0] _GEN_40 = 4'h0 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_0_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_41 = 4'h1 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_1_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_42 = 4'h2 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_2_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_43 = 4'h3 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_3_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_44 = 4'h4 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_4_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_45 = 4'h5 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_5_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_46 = 4'h6 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_6_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_47 = 4'h7 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_7_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_48 = 4'h8 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_8_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_49 = 4'h9 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_9_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_50 = 4'ha == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_10_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_51 = 4'hb == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_11_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_52 = 4'hc == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_12_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_53 = 4'hd == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_13_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_54 = 4'he == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_14_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_55 = 4'hf == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_15_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [33:0] _totalTx_memoryLength_T_1 = totalTx_memoryLength - 34'h40; // @[CScratchpad.scala 156:54]
  wire [33:0] _totalTx_memoryAddress_T_1 = totalTx_memoryAddress + 34'h40; // @[CScratchpad.scala 158:56]
  wire [1:0] _GEN_56 = isBelowLimit ? 2'h2 : mem_tx_state; // @[CScratchpad.scala 159:28 160:24 102:37]
  wire  _GEN_57 = _T_13 ? _GEN_8 : reqIdleBits_0; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_58 = _T_13 ? _GEN_9 : reqIdleBits_1; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_59 = _T_13 ? _GEN_10 : reqIdleBits_2; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_60 = _T_13 ? _GEN_11 : reqIdleBits_3; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_61 = _T_13 ? _GEN_12 : reqIdleBits_4; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_62 = _T_13 ? _GEN_13 : reqIdleBits_5; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_63 = _T_13 ? _GEN_14 : reqIdleBits_6; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_64 = _T_13 ? _GEN_15 : reqIdleBits_7; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_65 = _T_13 ? _GEN_16 : reqIdleBits_8; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_66 = _T_13 ? _GEN_17 : reqIdleBits_9; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_67 = _T_13 ? _GEN_18 : reqIdleBits_10; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_68 = _T_13 ? _GEN_19 : reqIdleBits_11; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_69 = _T_13 ? _GEN_20 : reqIdleBits_12; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_70 = _T_13 ? _GEN_21 : reqIdleBits_13; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_71 = _T_13 ? _GEN_22 : reqIdleBits_14; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_72 = _T_13 ? _GEN_23 : reqIdleBits_15; // @[CScratchpad.scala 152:28 110:36]
  wire [15:0] _GEN_89 = _T_13 ? _GEN_40 : req_cache_0_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_90 = _T_13 ? _GEN_41 : req_cache_1_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_91 = _T_13 ? _GEN_42 : req_cache_2_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_92 = _T_13 ? _GEN_43 : req_cache_3_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_93 = _T_13 ? _GEN_44 : req_cache_4_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_94 = _T_13 ? _GEN_45 : req_cache_5_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_95 = _T_13 ? _GEN_46 : req_cache_6_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_96 = _T_13 ? _GEN_47 : req_cache_7_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_97 = _T_13 ? _GEN_48 : req_cache_8_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_98 = _T_13 ? _GEN_49 : req_cache_9_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_99 = _T_13 ? _GEN_50 : req_cache_10_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_100 = _T_13 ? _GEN_51 : req_cache_11_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_101 = _T_13 ? _GEN_52 : req_cache_12_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_102 = _T_13 ? _GEN_53 : req_cache_13_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_103 = _T_13 ? _GEN_54 : req_cache_14_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_104 = _T_13 ? _GEN_55 : req_cache_15_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [1:0] _GEN_109 = reqIdleBits_0 & reqIdleBits_1 & reqIdleBits_2 & reqIdleBits_3 & reqIdleBits_4 & reqIdleBits_5 &
    reqIdleBits_6 & reqIdleBits_7 & reqIdleBits_8 & reqIdleBits_9 & reqIdleBits_10 & reqIdleBits_11 & reqIdleBits_12 &
    reqIdleBits_13 & reqIdleBits_14 & reqIdleBits_15 ? 2'h0 : mem_tx_state; // @[CScratchpad.scala 166:40 167:22 102:37]
  wire  _GEN_113 = 2'h1 == mem_tx_state ? _GEN_57 : reqIdleBits_0; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_114 = 2'h1 == mem_tx_state ? _GEN_58 : reqIdleBits_1; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_115 = 2'h1 == mem_tx_state ? _GEN_59 : reqIdleBits_2; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_116 = 2'h1 == mem_tx_state ? _GEN_60 : reqIdleBits_3; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_117 = 2'h1 == mem_tx_state ? _GEN_61 : reqIdleBits_4; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_118 = 2'h1 == mem_tx_state ? _GEN_62 : reqIdleBits_5; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_119 = 2'h1 == mem_tx_state ? _GEN_63 : reqIdleBits_6; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_120 = 2'h1 == mem_tx_state ? _GEN_64 : reqIdleBits_7; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_121 = 2'h1 == mem_tx_state ? _GEN_65 : reqIdleBits_8; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_122 = 2'h1 == mem_tx_state ? _GEN_66 : reqIdleBits_9; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_123 = 2'h1 == mem_tx_state ? _GEN_67 : reqIdleBits_10; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_124 = 2'h1 == mem_tx_state ? _GEN_68 : reqIdleBits_11; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_125 = 2'h1 == mem_tx_state ? _GEN_69 : reqIdleBits_12; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_126 = 2'h1 == mem_tx_state ? _GEN_70 : reqIdleBits_13; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_127 = 2'h1 == mem_tx_state ? _GEN_71 : reqIdleBits_14; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_128 = 2'h1 == mem_tx_state ? _GEN_72 : reqIdleBits_15; // @[CScratchpad.scala 138:24 110:36]
  wire [15:0] _GEN_145 = 2'h1 == mem_tx_state ? _GEN_89 : req_cache_0_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_146 = 2'h1 == mem_tx_state ? _GEN_90 : req_cache_1_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_147 = 2'h1 == mem_tx_state ? _GEN_91 : req_cache_2_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_148 = 2'h1 == mem_tx_state ? _GEN_92 : req_cache_3_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_149 = 2'h1 == mem_tx_state ? _GEN_93 : req_cache_4_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_150 = 2'h1 == mem_tx_state ? _GEN_94 : req_cache_5_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_151 = 2'h1 == mem_tx_state ? _GEN_95 : req_cache_6_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_152 = 2'h1 == mem_tx_state ? _GEN_96 : req_cache_7_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_153 = 2'h1 == mem_tx_state ? _GEN_97 : req_cache_8_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_154 = 2'h1 == mem_tx_state ? _GEN_98 : req_cache_9_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_155 = 2'h1 == mem_tx_state ? _GEN_99 : req_cache_10_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_156 = 2'h1 == mem_tx_state ? _GEN_100 : req_cache_11_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_157 = 2'h1 == mem_tx_state ? _GEN_101 : req_cache_12_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_158 = 2'h1 == mem_tx_state ? _GEN_102 : req_cache_13_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_159 = 2'h1 == mem_tx_state ? _GEN_103 : req_cache_14_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_160 = 2'h1 == mem_tx_state ? _GEN_104 : req_cache_15_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire  _GEN_171 = 2'h0 == mem_tx_state ? reqIdleBits_0 : _GEN_113; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_172 = 2'h0 == mem_tx_state ? reqIdleBits_1 : _GEN_114; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_173 = 2'h0 == mem_tx_state ? reqIdleBits_2 : _GEN_115; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_174 = 2'h0 == mem_tx_state ? reqIdleBits_3 : _GEN_116; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_175 = 2'h0 == mem_tx_state ? reqIdleBits_4 : _GEN_117; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_176 = 2'h0 == mem_tx_state ? reqIdleBits_5 : _GEN_118; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_177 = 2'h0 == mem_tx_state ? reqIdleBits_6 : _GEN_119; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_178 = 2'h0 == mem_tx_state ? reqIdleBits_7 : _GEN_120; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_179 = 2'h0 == mem_tx_state ? reqIdleBits_8 : _GEN_121; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_180 = 2'h0 == mem_tx_state ? reqIdleBits_9 : _GEN_122; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_181 = 2'h0 == mem_tx_state ? reqIdleBits_10 : _GEN_123; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_182 = 2'h0 == mem_tx_state ? reqIdleBits_11 : _GEN_124; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_183 = 2'h0 == mem_tx_state ? reqIdleBits_12 : _GEN_125; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_184 = 2'h0 == mem_tx_state ? reqIdleBits_13 : _GEN_126; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_185 = 2'h0 == mem_tx_state ? reqIdleBits_14 : _GEN_127; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_186 = 2'h0 == mem_tx_state ? reqIdleBits_15 : _GEN_128; // @[CScratchpad.scala 138:24 110:36]
  wire [15:0] _GEN_203 = 2'h0 == mem_tx_state ? req_cache_0_memoryLength : _GEN_145; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_204 = 2'h0 == mem_tx_state ? req_cache_1_memoryLength : _GEN_146; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_205 = 2'h0 == mem_tx_state ? req_cache_2_memoryLength : _GEN_147; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_206 = 2'h0 == mem_tx_state ? req_cache_3_memoryLength : _GEN_148; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_207 = 2'h0 == mem_tx_state ? req_cache_4_memoryLength : _GEN_149; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_208 = 2'h0 == mem_tx_state ? req_cache_5_memoryLength : _GEN_150; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_209 = 2'h0 == mem_tx_state ? req_cache_6_memoryLength : _GEN_151; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_210 = 2'h0 == mem_tx_state ? req_cache_7_memoryLength : _GEN_152; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_211 = 2'h0 == mem_tx_state ? req_cache_8_memoryLength : _GEN_153; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_212 = 2'h0 == mem_tx_state ? req_cache_9_memoryLength : _GEN_154; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_213 = 2'h0 == mem_tx_state ? req_cache_10_memoryLength : _GEN_155; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_214 = 2'h0 == mem_tx_state ? req_cache_11_memoryLength : _GEN_156; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_215 = 2'h0 == mem_tx_state ? req_cache_12_memoryLength : _GEN_157; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_216 = 2'h0 == mem_tx_state ? req_cache_13_memoryLength : _GEN_158; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_217 = 2'h0 == mem_tx_state ? req_cache_14_memoryLength : _GEN_159; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_218 = 2'h0 == mem_tx_state ? req_cache_15_memoryLength : _GEN_160; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_220 = 4'h1 == auto_mem_out_d_bits_source ? req_cache_1_memoryLength : req_cache_0_memoryLength; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_221 = 4'h2 == auto_mem_out_d_bits_source ? req_cache_2_memoryLength : _GEN_220; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_222 = 4'h3 == auto_mem_out_d_bits_source ? req_cache_3_memoryLength : _GEN_221; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_223 = 4'h4 == auto_mem_out_d_bits_source ? req_cache_4_memoryLength : _GEN_222; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_224 = 4'h5 == auto_mem_out_d_bits_source ? req_cache_5_memoryLength : _GEN_223; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_225 = 4'h6 == auto_mem_out_d_bits_source ? req_cache_6_memoryLength : _GEN_224; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_226 = 4'h7 == auto_mem_out_d_bits_source ? req_cache_7_memoryLength : _GEN_225; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_227 = 4'h8 == auto_mem_out_d_bits_source ? req_cache_8_memoryLength : _GEN_226; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_228 = 4'h9 == auto_mem_out_d_bits_source ? req_cache_9_memoryLength : _GEN_227; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_229 = 4'ha == auto_mem_out_d_bits_source ? req_cache_10_memoryLength : _GEN_228; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_230 = 4'hb == auto_mem_out_d_bits_source ? req_cache_11_memoryLength : _GEN_229; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_231 = 4'hc == auto_mem_out_d_bits_source ? req_cache_12_memoryLength : _GEN_230; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_232 = 4'hd == auto_mem_out_d_bits_source ? req_cache_13_memoryLength : _GEN_231; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_233 = 4'he == auto_mem_out_d_bits_source ? req_cache_14_memoryLength : _GEN_232; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_234 = 4'hf == auto_mem_out_d_bits_source ? req_cache_15_memoryLength : _GEN_233; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_235 = _GEN_234 >= 16'h40 ? 16'h40 : _GEN_234; // @[CScratchpad.scala 174:55 175:39 177:39]
  wire  mem_out_d_ready = loader_io_cache_block_in_ready; // @[Nodes.scala 1212:84 CScratchpad.scala 180:19]
  wire  _T_36 = mem_out_d_ready & auto_mem_out_d_valid; // @[Decoupled.scala 51:35]
  wire [15:0] _req_cache_memoryLength_T_2 = _GEN_234 - 16'h40; // @[CScratchpad.scala 210:72]
  wire  _GEN_445 = 4'h0 == auto_mem_out_d_bits_source | _GEN_171; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_446 = 4'h1 == auto_mem_out_d_bits_source | _GEN_172; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_447 = 4'h2 == auto_mem_out_d_bits_source | _GEN_173; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_448 = 4'h3 == auto_mem_out_d_bits_source | _GEN_174; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_449 = 4'h4 == auto_mem_out_d_bits_source | _GEN_175; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_450 = 4'h5 == auto_mem_out_d_bits_source | _GEN_176; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_451 = 4'h6 == auto_mem_out_d_bits_source | _GEN_177; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_452 = 4'h7 == auto_mem_out_d_bits_source | _GEN_178; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_453 = 4'h8 == auto_mem_out_d_bits_source | _GEN_179; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_454 = 4'h9 == auto_mem_out_d_bits_source | _GEN_180; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_455 = 4'ha == auto_mem_out_d_bits_source | _GEN_181; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_456 = 4'hb == auto_mem_out_d_bits_source | _GEN_182; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_457 = 4'hc == auto_mem_out_d_bits_source | _GEN_183; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_458 = 4'hd == auto_mem_out_d_bits_source | _GEN_184; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_459 = 4'he == auto_mem_out_d_bits_source | _GEN_185; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_460 = 4'hf == auto_mem_out_d_bits_source | _GEN_186; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_461 = _GEN_234 <= 16'h40 ? _GEN_445 : _GEN_171; // @[CScratchpad.scala 212:57]
  wire  _GEN_462 = _GEN_234 <= 16'h40 ? _GEN_446 : _GEN_172; // @[CScratchpad.scala 212:57]
  wire  _GEN_463 = _GEN_234 <= 16'h40 ? _GEN_447 : _GEN_173; // @[CScratchpad.scala 212:57]
  wire  _GEN_464 = _GEN_234 <= 16'h40 ? _GEN_448 : _GEN_174; // @[CScratchpad.scala 212:57]
  wire  _GEN_465 = _GEN_234 <= 16'h40 ? _GEN_449 : _GEN_175; // @[CScratchpad.scala 212:57]
  wire  _GEN_466 = _GEN_234 <= 16'h40 ? _GEN_450 : _GEN_176; // @[CScratchpad.scala 212:57]
  wire  _GEN_467 = _GEN_234 <= 16'h40 ? _GEN_451 : _GEN_177; // @[CScratchpad.scala 212:57]
  wire  _GEN_468 = _GEN_234 <= 16'h40 ? _GEN_452 : _GEN_178; // @[CScratchpad.scala 212:57]
  wire  _GEN_469 = _GEN_234 <= 16'h40 ? _GEN_453 : _GEN_179; // @[CScratchpad.scala 212:57]
  wire  _GEN_470 = _GEN_234 <= 16'h40 ? _GEN_454 : _GEN_180; // @[CScratchpad.scala 212:57]
  wire  _GEN_471 = _GEN_234 <= 16'h40 ? _GEN_455 : _GEN_181; // @[CScratchpad.scala 212:57]
  wire  _GEN_472 = _GEN_234 <= 16'h40 ? _GEN_456 : _GEN_182; // @[CScratchpad.scala 212:57]
  wire  _GEN_473 = _GEN_234 <= 16'h40 ? _GEN_457 : _GEN_183; // @[CScratchpad.scala 212:57]
  wire  _GEN_474 = _GEN_234 <= 16'h40 ? _GEN_458 : _GEN_184; // @[CScratchpad.scala 212:57]
  wire  _GEN_475 = _GEN_234 <= 16'h40 ? _GEN_459 : _GEN_185; // @[CScratchpad.scala 212:57]
  wire  _GEN_476 = _GEN_234 <= 16'h40 ? _GEN_460 : _GEN_186; // @[CScratchpad.scala 212:57]
  wire  _GEN_494 = _T_36 ? _GEN_461 : _GEN_171; // @[CScratchpad.scala 209:24]
  wire  _GEN_495 = _T_36 ? _GEN_462 : _GEN_172; // @[CScratchpad.scala 209:24]
  wire  _GEN_496 = _T_36 ? _GEN_463 : _GEN_173; // @[CScratchpad.scala 209:24]
  wire  _GEN_497 = _T_36 ? _GEN_464 : _GEN_174; // @[CScratchpad.scala 209:24]
  wire  _GEN_498 = _T_36 ? _GEN_465 : _GEN_175; // @[CScratchpad.scala 209:24]
  wire  _GEN_499 = _T_36 ? _GEN_466 : _GEN_176; // @[CScratchpad.scala 209:24]
  wire  _GEN_500 = _T_36 ? _GEN_467 : _GEN_177; // @[CScratchpad.scala 209:24]
  wire  _GEN_501 = _T_36 ? _GEN_468 : _GEN_178; // @[CScratchpad.scala 209:24]
  wire  _GEN_502 = _T_36 ? _GEN_469 : _GEN_179; // @[CScratchpad.scala 209:24]
  wire  _GEN_503 = _T_36 ? _GEN_470 : _GEN_180; // @[CScratchpad.scala 209:24]
  wire  _GEN_504 = _T_36 ? _GEN_471 : _GEN_181; // @[CScratchpad.scala 209:24]
  wire  _GEN_505 = _T_36 ? _GEN_472 : _GEN_182; // @[CScratchpad.scala 209:24]
  wire  _GEN_506 = _T_36 ? _GEN_473 : _GEN_183; // @[CScratchpad.scala 209:24]
  wire  _GEN_507 = _T_36 ? _GEN_474 : _GEN_184; // @[CScratchpad.scala 209:24]
  wire  _GEN_508 = _T_36 ? _GEN_475 : _GEN_185; // @[CScratchpad.scala 209:24]
  wire  _GEN_509 = _T_36 ? _GEN_476 : _GEN_186; // @[CScratchpad.scala 209:24]
  CScratchpadPackedSubwordLoader_2 loader ( // @[CScratchpad.scala 94:30]
    .clock(loader_clock),
    .reset(loader_reset),
    .io_cache_block_in_ready(loader_io_cache_block_in_ready),
    .io_cache_block_in_valid(loader_io_cache_block_in_valid),
    .io_cache_block_in_bits_len(loader_io_cache_block_in_bits_len),
    .io_sp_write_out_valid(loader_io_sp_write_out_valid)
  );
  assign auto_mem_out_a_valid = 2'h0 == mem_tx_state ? mem_tx_state == 2'h1 : _GEN_112; // @[CScratchpad.scala 136:19 138:24]
  assign auto_mem_out_a_bits_size = txEmitLengthLg[2:0]; // @[Edges.scala 447:17 450:15]
  assign auto_mem_out_a_bits_source = reqIdleBits_0 ? 4'h0 : _reqChosen_T_13; // @[Mux.scala 47:70]
  assign auto_mem_out_a_bits_address = totalTx_memoryAddress; // @[Edges.scala 447:17 452:15]
  assign auto_mem_out_a_bits_mask = {x1_a_bits_a_mask_hi,x1_a_bits_a_mask_lo}; // @[Cat.scala 33:92]
  assign auto_mem_out_d_ready = loader_io_cache_block_in_ready; // @[Nodes.scala 1212:84 CScratchpad.scala 180:19]
  assign loader_clock = clock;
  assign loader_reset = reset;
  assign loader_io_cache_block_in_valid = auto_mem_out_d_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign loader_io_cache_block_in_bits_len = _GEN_235[6:0];
  always @(posedge clock) begin
    if (reset) begin // @[CScratchpad.scala 102:37]
      mem_tx_state <= 2'h0; // @[CScratchpad.scala 102:37]
    end else if (!(2'h0 == mem_tx_state)) begin // @[CScratchpad.scala 138:24]
      if (2'h1 == mem_tx_state) begin // @[CScratchpad.scala 138:24]
        if (_T_13) begin // @[CScratchpad.scala 152:28]
          mem_tx_state <= _GEN_56;
        end
      end else if (2'h2 == mem_tx_state) begin // @[CScratchpad.scala 138:24]
        mem_tx_state <= _GEN_109;
      end
    end
    reqIdleBits_0 <= reset | _GEN_494; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_1 <= reset | _GEN_495; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_2 <= reset | _GEN_496; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_3 <= reset | _GEN_497; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_4 <= reset | _GEN_498; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_5 <= reset | _GEN_499; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_6 <= reset | _GEN_500; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_7 <= reset | _GEN_501; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_8 <= reset | _GEN_502; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_9 <= reset | _GEN_503; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_10 <= reset | _GEN_504; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_11 <= reset | _GEN_505; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_12 <= reset | _GEN_506; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_13 <= reset | _GEN_507; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_14 <= reset | _GEN_508; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_15 <= reset | _GEN_509; // @[CScratchpad.scala 110:{36,36}]
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h0 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_0_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_0_memoryLength <= _GEN_203;
      end
    end else begin
      req_cache_0_memoryLength <= _GEN_203;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h1 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_1_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_1_memoryLength <= _GEN_204;
      end
    end else begin
      req_cache_1_memoryLength <= _GEN_204;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h2 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_2_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_2_memoryLength <= _GEN_205;
      end
    end else begin
      req_cache_2_memoryLength <= _GEN_205;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h3 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_3_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_3_memoryLength <= _GEN_206;
      end
    end else begin
      req_cache_3_memoryLength <= _GEN_206;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h4 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_4_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_4_memoryLength <= _GEN_207;
      end
    end else begin
      req_cache_4_memoryLength <= _GEN_207;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h5 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_5_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_5_memoryLength <= _GEN_208;
      end
    end else begin
      req_cache_5_memoryLength <= _GEN_208;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h6 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_6_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_6_memoryLength <= _GEN_209;
      end
    end else begin
      req_cache_6_memoryLength <= _GEN_209;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h7 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_7_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_7_memoryLength <= _GEN_210;
      end
    end else begin
      req_cache_7_memoryLength <= _GEN_210;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h8 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_8_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_8_memoryLength <= _GEN_211;
      end
    end else begin
      req_cache_8_memoryLength <= _GEN_211;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h9 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_9_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_9_memoryLength <= _GEN_212;
      end
    end else begin
      req_cache_9_memoryLength <= _GEN_212;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'ha == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_10_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_10_memoryLength <= _GEN_213;
      end
    end else begin
      req_cache_10_memoryLength <= _GEN_213;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'hb == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_11_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_11_memoryLength <= _GEN_214;
      end
    end else begin
      req_cache_11_memoryLength <= _GEN_214;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'hc == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_12_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_12_memoryLength <= _GEN_215;
      end
    end else begin
      req_cache_12_memoryLength <= _GEN_215;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'hd == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_13_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_13_memoryLength <= _GEN_216;
      end
    end else begin
      req_cache_13_memoryLength <= _GEN_216;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'he == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_14_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_14_memoryLength <= _GEN_217;
      end
    end else begin
      req_cache_14_memoryLength <= _GEN_217;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'hf == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_15_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_15_memoryLength <= _GEN_218;
      end
    end else begin
      req_cache_15_memoryLength <= _GEN_218;
    end
    if (!(2'h0 == mem_tx_state)) begin // @[CScratchpad.scala 138:24]
      if (2'h1 == mem_tx_state) begin // @[CScratchpad.scala 138:24]
        if (_T_13) begin // @[CScratchpad.scala 152:28]
          totalTx_memoryAddress <= _totalTx_memoryAddress_T_1; // @[CScratchpad.scala 158:31]
        end
      end
    end
    if (!(2'h0 == mem_tx_state)) begin // @[CScratchpad.scala 138:24]
      if (2'h1 == mem_tx_state) begin // @[CScratchpad.scala 138:24]
        if (_T_13) begin // @[CScratchpad.scala 152:28]
          totalTx_memoryLength <= _totalTx_memoryLength_T_1; // @[CScratchpad.scala 156:30]
        end
      end
    end
  end
endmodule
module CScratchpadPackedSubwordLoader_3(
  input        clock,
  input        reset,
  output       io_cache_block_in_ready,
  input        io_cache_block_in_valid,
  input  [6:0] io_cache_block_in_bits_len,
  output       io_sp_write_out_valid
);
  reg [6:0] lenRemainingFromReq; // @[CScratchpadPackedSubwordLoader.scala 18:32]
  reg  state; // @[CScratchpadPackedSubwordLoader.scala 21:22]
  wire  _io_cache_block_in_ready_T = ~state; // @[CScratchpadPackedSubwordLoader.scala 22:36]
  wire  _T_1 = io_cache_block_in_ready & io_cache_block_in_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_0 = _T_1 | state; // @[CScratchpadPackedSubwordLoader.scala 34:36 35:15 21:22]
  wire [6:0] _lenRemainingFromReq_T_1 = lenRemainingFromReq - 7'h20; // @[CScratchpadPackedSubwordLoader.scala 53:54]
  wire  _GEN_6 = lenRemainingFromReq == 7'h20 ? 1'h0 : state; // @[CScratchpadPackedSubwordLoader.scala 54:60 55:19 21:22]
  assign io_cache_block_in_ready = ~state; // @[CScratchpadPackedSubwordLoader.scala 22:36]
  assign io_sp_write_out_valid = _io_cache_block_in_ready_T ? 1'h0 : state; // @[CScratchpadPackedSubwordLoader.scala 32:17 24:25]
  always @(posedge clock) begin
    if (_io_cache_block_in_ready_T) begin // @[CScratchpadPackedSubwordLoader.scala 32:17]
      if (_T_1) begin // @[CScratchpadPackedSubwordLoader.scala 34:36]
        lenRemainingFromReq <= io_cache_block_in_bits_len; // @[CScratchpadPackedSubwordLoader.scala 38:29]
      end
    end else if (state) begin // @[CScratchpadPackedSubwordLoader.scala 32:17]
      if (io_sp_write_out_valid) begin // @[CScratchpadPackedSubwordLoader.scala 48:34]
        lenRemainingFromReq <= _lenRemainingFromReq_T_1;
      end
    end
    if (reset) begin // @[CScratchpadPackedSubwordLoader.scala 21:22]
      state <= 1'h0; // @[CScratchpadPackedSubwordLoader.scala 21:22]
    end else if (_io_cache_block_in_ready_T) begin // @[CScratchpadPackedSubwordLoader.scala 32:17]
      state <= _GEN_0;
    end else if (state) begin // @[CScratchpadPackedSubwordLoader.scala 32:17]
      if (io_sp_write_out_valid) begin // @[CScratchpadPackedSubwordLoader.scala 48:34]
        state <= _GEN_6;
      end
    end
  end
endmodule
module CScratchpad_3(
  input         clock,
  input         reset,
  input         auto_mem_out_a_ready,
  output        auto_mem_out_a_valid,
  output [2:0]  auto_mem_out_a_bits_size,
  output [3:0]  auto_mem_out_a_bits_source,
  output [33:0] auto_mem_out_a_bits_address,
  output [63:0] auto_mem_out_a_bits_mask,
  output        auto_mem_out_d_ready,
  input         auto_mem_out_d_valid,
  input  [3:0]  auto_mem_out_d_bits_source
);
  wire  loader_clock; // @[CScratchpad.scala 94:30]
  wire  loader_reset; // @[CScratchpad.scala 94:30]
  wire  loader_io_cache_block_in_ready; // @[CScratchpad.scala 94:30]
  wire  loader_io_cache_block_in_valid; // @[CScratchpad.scala 94:30]
  wire [6:0] loader_io_cache_block_in_bits_len; // @[CScratchpad.scala 94:30]
  wire  loader_io_sp_write_out_valid; // @[CScratchpad.scala 94:30]
  reg [1:0] mem_tx_state; // @[CScratchpad.scala 102:37]
  reg  reqIdleBits_0; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_1; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_2; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_3; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_4; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_5; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_6; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_7; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_8; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_9; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_10; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_11; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_12; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_13; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_14; // @[CScratchpad.scala 110:36]
  reg  reqIdleBits_15; // @[CScratchpad.scala 110:36]
  wire  reqAvailable = reqIdleBits_0 | reqIdleBits_1 | reqIdleBits_2 | reqIdleBits_3 | reqIdleBits_4 | reqIdleBits_5 |
    reqIdleBits_6 | reqIdleBits_7 | reqIdleBits_8 | reqIdleBits_9 | reqIdleBits_10 | reqIdleBits_11 | reqIdleBits_12 |
    reqIdleBits_13 | reqIdleBits_14 | reqIdleBits_15; // @[CScratchpad.scala 111:51]
  wire [3:0] _reqChosen_T = reqIdleBits_14 ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_1 = reqIdleBits_13 ? 4'hd : _reqChosen_T; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_2 = reqIdleBits_12 ? 4'hc : _reqChosen_T_1; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_3 = reqIdleBits_11 ? 4'hb : _reqChosen_T_2; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_4 = reqIdleBits_10 ? 4'ha : _reqChosen_T_3; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_5 = reqIdleBits_9 ? 4'h9 : _reqChosen_T_4; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_6 = reqIdleBits_8 ? 4'h8 : _reqChosen_T_5; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_7 = reqIdleBits_7 ? 4'h7 : _reqChosen_T_6; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_8 = reqIdleBits_6 ? 4'h6 : _reqChosen_T_7; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_9 = reqIdleBits_5 ? 4'h5 : _reqChosen_T_8; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_10 = reqIdleBits_4 ? 4'h4 : _reqChosen_T_9; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_11 = reqIdleBits_3 ? 4'h3 : _reqChosen_T_10; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_12 = reqIdleBits_2 ? 4'h2 : _reqChosen_T_11; // @[Mux.scala 47:70]
  wire [3:0] _reqChosen_T_13 = reqIdleBits_1 ? 4'h1 : _reqChosen_T_12; // @[Mux.scala 47:70]
  wire [3:0] reqChosen = reqIdleBits_0 ? 4'h0 : _reqChosen_T_13; // @[Mux.scala 47:70]
  reg [15:0] req_cache_0_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_1_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_2_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_3_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_4_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_5_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_6_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_7_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_8_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_9_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_10_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_11_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_12_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_13_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_14_memoryLength; // @[CScratchpad.scala 114:30]
  reg [15:0] req_cache_15_memoryLength; // @[CScratchpad.scala 114:30]
  reg [33:0] totalTx_memoryAddress; // @[CScratchpad.scala 124:28]
  reg [33:0] totalTx_memoryLength; // @[CScratchpad.scala 124:28]
  wire  isBelowLimit = totalTx_memoryLength <= 34'h40; // @[CScratchpad.scala 149:47]
  wire [1:0] txEmitLengthLg_hi = totalTx_memoryLength[33:32]; // @[OneHot.scala 30:18]
  wire  _txEmitLengthLg_T = |txEmitLengthLg_hi; // @[OneHot.scala 32:14]
  wire [31:0] txEmitLengthLg_lo = totalTx_memoryLength[31:0]; // @[OneHot.scala 31:18]
  wire [31:0] _GEN_569 = {{30'd0}, txEmitLengthLg_hi}; // @[OneHot.scala 32:28]
  wire [31:0] _txEmitLengthLg_T_1 = _GEN_569 | txEmitLengthLg_lo; // @[OneHot.scala 32:28]
  wire [15:0] txEmitLengthLg_hi_1 = _txEmitLengthLg_T_1[31:16]; // @[OneHot.scala 30:18]
  wire  _txEmitLengthLg_T_2 = |txEmitLengthLg_hi_1; // @[OneHot.scala 32:14]
  wire [15:0] txEmitLengthLg_lo_1 = _txEmitLengthLg_T_1[15:0]; // @[OneHot.scala 31:18]
  wire [15:0] _txEmitLengthLg_T_3 = txEmitLengthLg_hi_1 | txEmitLengthLg_lo_1; // @[OneHot.scala 32:28]
  wire [7:0] txEmitLengthLg_hi_2 = _txEmitLengthLg_T_3[15:8]; // @[OneHot.scala 30:18]
  wire  _txEmitLengthLg_T_4 = |txEmitLengthLg_hi_2; // @[OneHot.scala 32:14]
  wire [7:0] txEmitLengthLg_lo_2 = _txEmitLengthLg_T_3[7:0]; // @[OneHot.scala 31:18]
  wire [7:0] _txEmitLengthLg_T_5 = txEmitLengthLg_hi_2 | txEmitLengthLg_lo_2; // @[OneHot.scala 32:28]
  wire [3:0] txEmitLengthLg_hi_3 = _txEmitLengthLg_T_5[7:4]; // @[OneHot.scala 30:18]
  wire  _txEmitLengthLg_T_6 = |txEmitLengthLg_hi_3; // @[OneHot.scala 32:14]
  wire [3:0] txEmitLengthLg_lo_3 = _txEmitLengthLg_T_5[3:0]; // @[OneHot.scala 31:18]
  wire [3:0] _txEmitLengthLg_T_7 = txEmitLengthLg_hi_3 | txEmitLengthLg_lo_3; // @[OneHot.scala 32:28]
  wire [1:0] txEmitLengthLg_hi_4 = _txEmitLengthLg_T_7[3:2]; // @[OneHot.scala 30:18]
  wire  _txEmitLengthLg_T_8 = |txEmitLengthLg_hi_4; // @[OneHot.scala 32:14]
  wire [1:0] txEmitLengthLg_lo_4 = _txEmitLengthLg_T_7[1:0]; // @[OneHot.scala 31:18]
  wire [1:0] _txEmitLengthLg_T_9 = txEmitLengthLg_hi_4 | txEmitLengthLg_lo_4; // @[OneHot.scala 32:28]
  wire [5:0] _txEmitLengthLg_T_15 = {_txEmitLengthLg_T,_txEmitLengthLg_T_2,_txEmitLengthLg_T_4,_txEmitLengthLg_T_6,
    _txEmitLengthLg_T_8,_txEmitLengthLg_T_9[1]}; // @[Cat.scala 33:92]
  wire [5:0] _txEmitLengthLg_T_16 = isBelowLimit ? _txEmitLengthLg_T_15 : 6'h6; // @[CScratchpad.scala 150:28]
  wire [5:0] _GEN_111 = 2'h1 == mem_tx_state ? _txEmitLengthLg_T_16 : 6'h0; // @[CScratchpad.scala 131:18 138:24 150:22]
  wire [5:0] _GEN_169 = 2'h0 == mem_tx_state ? 6'h0 : _GEN_111; // @[CScratchpad.scala 131:18 138:24]
  wire [3:0] txEmitLengthLg = _GEN_169[3:0]; // @[CScratchpad.scala 130:36]
  wire [5:0] _x1_a_bits_a_mask_sizeOH_T = {{2'd0}, txEmitLengthLg}; // @[Misc.scala 201:34]
  wire [2:0] x1_a_bits_a_mask_sizeOH_shiftAmount = _x1_a_bits_a_mask_sizeOH_T[2:0]; // @[OneHot.scala 63:49]
  wire [7:0] _x1_a_bits_a_mask_sizeOH_T_1 = 8'h1 << x1_a_bits_a_mask_sizeOH_shiftAmount; // @[OneHot.scala 64:12]
  wire [5:0] x1_a_bits_a_mask_sizeOH = _x1_a_bits_a_mask_sizeOH_T_1[5:0] | 6'h1; // @[Misc.scala 201:81]
  wire  _x1_a_bits_a_mask_T = txEmitLengthLg >= 4'h6; // @[Misc.scala 205:21]
  wire  x1_a_bits_a_mask_size = x1_a_bits_a_mask_sizeOH[5]; // @[Misc.scala 208:26]
  wire  x1_a_bits_a_mask_bit = totalTx_memoryAddress[5]; // @[Misc.scala 209:26]
  wire  x1_a_bits_a_mask_nbit = ~x1_a_bits_a_mask_bit; // @[Misc.scala 210:20]
  wire  x1_a_bits_a_mask_acc = _x1_a_bits_a_mask_T | x1_a_bits_a_mask_size & x1_a_bits_a_mask_nbit; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_acc_1 = _x1_a_bits_a_mask_T | x1_a_bits_a_mask_size & x1_a_bits_a_mask_bit; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_size_1 = x1_a_bits_a_mask_sizeOH[4]; // @[Misc.scala 208:26]
  wire  x1_a_bits_a_mask_bit_1 = totalTx_memoryAddress[4]; // @[Misc.scala 209:26]
  wire  x1_a_bits_a_mask_nbit_1 = ~x1_a_bits_a_mask_bit_1; // @[Misc.scala 210:20]
  wire  x1_a_bits_a_mask_eq_2 = x1_a_bits_a_mask_nbit & x1_a_bits_a_mask_nbit_1; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_2 = x1_a_bits_a_mask_acc | x1_a_bits_a_mask_size_1 & x1_a_bits_a_mask_eq_2; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_3 = x1_a_bits_a_mask_nbit & x1_a_bits_a_mask_bit_1; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_3 = x1_a_bits_a_mask_acc | x1_a_bits_a_mask_size_1 & x1_a_bits_a_mask_eq_3; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_4 = x1_a_bits_a_mask_bit & x1_a_bits_a_mask_nbit_1; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_4 = x1_a_bits_a_mask_acc_1 | x1_a_bits_a_mask_size_1 & x1_a_bits_a_mask_eq_4; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_5 = x1_a_bits_a_mask_bit & x1_a_bits_a_mask_bit_1; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_5 = x1_a_bits_a_mask_acc_1 | x1_a_bits_a_mask_size_1 & x1_a_bits_a_mask_eq_5; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_size_2 = x1_a_bits_a_mask_sizeOH[3]; // @[Misc.scala 208:26]
  wire  x1_a_bits_a_mask_bit_2 = totalTx_memoryAddress[3]; // @[Misc.scala 209:26]
  wire  x1_a_bits_a_mask_nbit_2 = ~x1_a_bits_a_mask_bit_2; // @[Misc.scala 210:20]
  wire  x1_a_bits_a_mask_eq_6 = x1_a_bits_a_mask_eq_2 & x1_a_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_6 = x1_a_bits_a_mask_acc_2 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_6; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_7 = x1_a_bits_a_mask_eq_2 & x1_a_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_7 = x1_a_bits_a_mask_acc_2 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_7; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_8 = x1_a_bits_a_mask_eq_3 & x1_a_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_8 = x1_a_bits_a_mask_acc_3 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_8; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_9 = x1_a_bits_a_mask_eq_3 & x1_a_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_9 = x1_a_bits_a_mask_acc_3 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_9; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_10 = x1_a_bits_a_mask_eq_4 & x1_a_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_10 = x1_a_bits_a_mask_acc_4 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_10; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_11 = x1_a_bits_a_mask_eq_4 & x1_a_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_11 = x1_a_bits_a_mask_acc_4 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_11; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_12 = x1_a_bits_a_mask_eq_5 & x1_a_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_12 = x1_a_bits_a_mask_acc_5 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_12; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_13 = x1_a_bits_a_mask_eq_5 & x1_a_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_13 = x1_a_bits_a_mask_acc_5 | x1_a_bits_a_mask_size_2 & x1_a_bits_a_mask_eq_13; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_size_3 = x1_a_bits_a_mask_sizeOH[2]; // @[Misc.scala 208:26]
  wire  x1_a_bits_a_mask_bit_3 = totalTx_memoryAddress[2]; // @[Misc.scala 209:26]
  wire  x1_a_bits_a_mask_nbit_3 = ~x1_a_bits_a_mask_bit_3; // @[Misc.scala 210:20]
  wire  x1_a_bits_a_mask_eq_14 = x1_a_bits_a_mask_eq_6 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_14 = x1_a_bits_a_mask_acc_6 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_14; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_15 = x1_a_bits_a_mask_eq_6 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_15 = x1_a_bits_a_mask_acc_6 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_15; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_16 = x1_a_bits_a_mask_eq_7 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_16 = x1_a_bits_a_mask_acc_7 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_16; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_17 = x1_a_bits_a_mask_eq_7 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_17 = x1_a_bits_a_mask_acc_7 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_17; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_18 = x1_a_bits_a_mask_eq_8 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_18 = x1_a_bits_a_mask_acc_8 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_18; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_19 = x1_a_bits_a_mask_eq_8 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_19 = x1_a_bits_a_mask_acc_8 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_19; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_20 = x1_a_bits_a_mask_eq_9 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_20 = x1_a_bits_a_mask_acc_9 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_20; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_21 = x1_a_bits_a_mask_eq_9 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_21 = x1_a_bits_a_mask_acc_9 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_21; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_22 = x1_a_bits_a_mask_eq_10 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_22 = x1_a_bits_a_mask_acc_10 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_22; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_23 = x1_a_bits_a_mask_eq_10 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_23 = x1_a_bits_a_mask_acc_10 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_23; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_24 = x1_a_bits_a_mask_eq_11 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_24 = x1_a_bits_a_mask_acc_11 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_24; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_25 = x1_a_bits_a_mask_eq_11 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_25 = x1_a_bits_a_mask_acc_11 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_25; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_26 = x1_a_bits_a_mask_eq_12 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_26 = x1_a_bits_a_mask_acc_12 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_26; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_27 = x1_a_bits_a_mask_eq_12 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_27 = x1_a_bits_a_mask_acc_12 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_27; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_28 = x1_a_bits_a_mask_eq_13 & x1_a_bits_a_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_28 = x1_a_bits_a_mask_acc_13 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_28; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_29 = x1_a_bits_a_mask_eq_13 & x1_a_bits_a_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_29 = x1_a_bits_a_mask_acc_13 | x1_a_bits_a_mask_size_3 & x1_a_bits_a_mask_eq_29; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_size_4 = x1_a_bits_a_mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  x1_a_bits_a_mask_bit_4 = totalTx_memoryAddress[1]; // @[Misc.scala 209:26]
  wire  x1_a_bits_a_mask_nbit_4 = ~x1_a_bits_a_mask_bit_4; // @[Misc.scala 210:20]
  wire  x1_a_bits_a_mask_eq_30 = x1_a_bits_a_mask_eq_14 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_30 = x1_a_bits_a_mask_acc_14 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_30; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_31 = x1_a_bits_a_mask_eq_14 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_31 = x1_a_bits_a_mask_acc_14 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_31; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_32 = x1_a_bits_a_mask_eq_15 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_32 = x1_a_bits_a_mask_acc_15 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_32; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_33 = x1_a_bits_a_mask_eq_15 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_33 = x1_a_bits_a_mask_acc_15 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_33; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_34 = x1_a_bits_a_mask_eq_16 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_34 = x1_a_bits_a_mask_acc_16 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_34; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_35 = x1_a_bits_a_mask_eq_16 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_35 = x1_a_bits_a_mask_acc_16 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_35; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_36 = x1_a_bits_a_mask_eq_17 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_36 = x1_a_bits_a_mask_acc_17 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_36; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_37 = x1_a_bits_a_mask_eq_17 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_37 = x1_a_bits_a_mask_acc_17 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_37; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_38 = x1_a_bits_a_mask_eq_18 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_38 = x1_a_bits_a_mask_acc_18 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_38; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_39 = x1_a_bits_a_mask_eq_18 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_39 = x1_a_bits_a_mask_acc_18 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_39; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_40 = x1_a_bits_a_mask_eq_19 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_40 = x1_a_bits_a_mask_acc_19 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_40; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_41 = x1_a_bits_a_mask_eq_19 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_41 = x1_a_bits_a_mask_acc_19 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_41; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_42 = x1_a_bits_a_mask_eq_20 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_42 = x1_a_bits_a_mask_acc_20 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_42; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_43 = x1_a_bits_a_mask_eq_20 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_43 = x1_a_bits_a_mask_acc_20 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_43; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_44 = x1_a_bits_a_mask_eq_21 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_44 = x1_a_bits_a_mask_acc_21 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_44; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_45 = x1_a_bits_a_mask_eq_21 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_45 = x1_a_bits_a_mask_acc_21 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_45; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_46 = x1_a_bits_a_mask_eq_22 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_46 = x1_a_bits_a_mask_acc_22 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_46; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_47 = x1_a_bits_a_mask_eq_22 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_47 = x1_a_bits_a_mask_acc_22 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_47; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_48 = x1_a_bits_a_mask_eq_23 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_48 = x1_a_bits_a_mask_acc_23 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_48; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_49 = x1_a_bits_a_mask_eq_23 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_49 = x1_a_bits_a_mask_acc_23 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_49; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_50 = x1_a_bits_a_mask_eq_24 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_50 = x1_a_bits_a_mask_acc_24 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_50; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_51 = x1_a_bits_a_mask_eq_24 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_51 = x1_a_bits_a_mask_acc_24 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_51; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_52 = x1_a_bits_a_mask_eq_25 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_52 = x1_a_bits_a_mask_acc_25 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_52; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_53 = x1_a_bits_a_mask_eq_25 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_53 = x1_a_bits_a_mask_acc_25 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_53; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_54 = x1_a_bits_a_mask_eq_26 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_54 = x1_a_bits_a_mask_acc_26 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_54; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_55 = x1_a_bits_a_mask_eq_26 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_55 = x1_a_bits_a_mask_acc_26 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_55; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_56 = x1_a_bits_a_mask_eq_27 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_56 = x1_a_bits_a_mask_acc_27 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_56; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_57 = x1_a_bits_a_mask_eq_27 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_57 = x1_a_bits_a_mask_acc_27 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_57; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_58 = x1_a_bits_a_mask_eq_28 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_58 = x1_a_bits_a_mask_acc_28 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_58; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_59 = x1_a_bits_a_mask_eq_28 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_59 = x1_a_bits_a_mask_acc_28 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_59; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_60 = x1_a_bits_a_mask_eq_29 & x1_a_bits_a_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_60 = x1_a_bits_a_mask_acc_29 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_60; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_61 = x1_a_bits_a_mask_eq_29 & x1_a_bits_a_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_61 = x1_a_bits_a_mask_acc_29 | x1_a_bits_a_mask_size_4 & x1_a_bits_a_mask_eq_61; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_size_5 = x1_a_bits_a_mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  x1_a_bits_a_mask_bit_5 = totalTx_memoryAddress[0]; // @[Misc.scala 209:26]
  wire  x1_a_bits_a_mask_nbit_5 = ~x1_a_bits_a_mask_bit_5; // @[Misc.scala 210:20]
  wire  x1_a_bits_a_mask_eq_62 = x1_a_bits_a_mask_eq_30 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_62 = x1_a_bits_a_mask_acc_30 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_62; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_63 = x1_a_bits_a_mask_eq_30 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_63 = x1_a_bits_a_mask_acc_30 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_63; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_64 = x1_a_bits_a_mask_eq_31 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_64 = x1_a_bits_a_mask_acc_31 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_64; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_65 = x1_a_bits_a_mask_eq_31 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_65 = x1_a_bits_a_mask_acc_31 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_65; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_66 = x1_a_bits_a_mask_eq_32 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_66 = x1_a_bits_a_mask_acc_32 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_66; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_67 = x1_a_bits_a_mask_eq_32 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_67 = x1_a_bits_a_mask_acc_32 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_67; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_68 = x1_a_bits_a_mask_eq_33 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_68 = x1_a_bits_a_mask_acc_33 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_68; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_69 = x1_a_bits_a_mask_eq_33 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_69 = x1_a_bits_a_mask_acc_33 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_69; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_70 = x1_a_bits_a_mask_eq_34 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_70 = x1_a_bits_a_mask_acc_34 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_70; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_71 = x1_a_bits_a_mask_eq_34 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_71 = x1_a_bits_a_mask_acc_34 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_71; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_72 = x1_a_bits_a_mask_eq_35 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_72 = x1_a_bits_a_mask_acc_35 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_72; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_73 = x1_a_bits_a_mask_eq_35 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_73 = x1_a_bits_a_mask_acc_35 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_73; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_74 = x1_a_bits_a_mask_eq_36 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_74 = x1_a_bits_a_mask_acc_36 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_74; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_75 = x1_a_bits_a_mask_eq_36 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_75 = x1_a_bits_a_mask_acc_36 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_75; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_76 = x1_a_bits_a_mask_eq_37 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_76 = x1_a_bits_a_mask_acc_37 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_76; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_77 = x1_a_bits_a_mask_eq_37 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_77 = x1_a_bits_a_mask_acc_37 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_77; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_78 = x1_a_bits_a_mask_eq_38 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_78 = x1_a_bits_a_mask_acc_38 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_78; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_79 = x1_a_bits_a_mask_eq_38 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_79 = x1_a_bits_a_mask_acc_38 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_79; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_80 = x1_a_bits_a_mask_eq_39 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_80 = x1_a_bits_a_mask_acc_39 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_80; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_81 = x1_a_bits_a_mask_eq_39 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_81 = x1_a_bits_a_mask_acc_39 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_81; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_82 = x1_a_bits_a_mask_eq_40 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_82 = x1_a_bits_a_mask_acc_40 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_82; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_83 = x1_a_bits_a_mask_eq_40 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_83 = x1_a_bits_a_mask_acc_40 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_83; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_84 = x1_a_bits_a_mask_eq_41 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_84 = x1_a_bits_a_mask_acc_41 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_84; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_85 = x1_a_bits_a_mask_eq_41 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_85 = x1_a_bits_a_mask_acc_41 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_85; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_86 = x1_a_bits_a_mask_eq_42 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_86 = x1_a_bits_a_mask_acc_42 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_86; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_87 = x1_a_bits_a_mask_eq_42 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_87 = x1_a_bits_a_mask_acc_42 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_87; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_88 = x1_a_bits_a_mask_eq_43 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_88 = x1_a_bits_a_mask_acc_43 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_88; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_89 = x1_a_bits_a_mask_eq_43 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_89 = x1_a_bits_a_mask_acc_43 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_89; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_90 = x1_a_bits_a_mask_eq_44 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_90 = x1_a_bits_a_mask_acc_44 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_90; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_91 = x1_a_bits_a_mask_eq_44 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_91 = x1_a_bits_a_mask_acc_44 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_91; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_92 = x1_a_bits_a_mask_eq_45 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_92 = x1_a_bits_a_mask_acc_45 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_92; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_93 = x1_a_bits_a_mask_eq_45 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_93 = x1_a_bits_a_mask_acc_45 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_93; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_94 = x1_a_bits_a_mask_eq_46 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_94 = x1_a_bits_a_mask_acc_46 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_94; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_95 = x1_a_bits_a_mask_eq_46 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_95 = x1_a_bits_a_mask_acc_46 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_95; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_96 = x1_a_bits_a_mask_eq_47 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_96 = x1_a_bits_a_mask_acc_47 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_96; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_97 = x1_a_bits_a_mask_eq_47 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_97 = x1_a_bits_a_mask_acc_47 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_97; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_98 = x1_a_bits_a_mask_eq_48 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_98 = x1_a_bits_a_mask_acc_48 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_98; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_99 = x1_a_bits_a_mask_eq_48 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_99 = x1_a_bits_a_mask_acc_48 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_99; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_100 = x1_a_bits_a_mask_eq_49 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_100 = x1_a_bits_a_mask_acc_49 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_100; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_101 = x1_a_bits_a_mask_eq_49 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_101 = x1_a_bits_a_mask_acc_49 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_101; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_102 = x1_a_bits_a_mask_eq_50 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_102 = x1_a_bits_a_mask_acc_50 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_102; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_103 = x1_a_bits_a_mask_eq_50 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_103 = x1_a_bits_a_mask_acc_50 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_103; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_104 = x1_a_bits_a_mask_eq_51 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_104 = x1_a_bits_a_mask_acc_51 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_104; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_105 = x1_a_bits_a_mask_eq_51 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_105 = x1_a_bits_a_mask_acc_51 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_105; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_106 = x1_a_bits_a_mask_eq_52 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_106 = x1_a_bits_a_mask_acc_52 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_106; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_107 = x1_a_bits_a_mask_eq_52 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_107 = x1_a_bits_a_mask_acc_52 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_107; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_108 = x1_a_bits_a_mask_eq_53 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_108 = x1_a_bits_a_mask_acc_53 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_108; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_109 = x1_a_bits_a_mask_eq_53 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_109 = x1_a_bits_a_mask_acc_53 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_109; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_110 = x1_a_bits_a_mask_eq_54 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_110 = x1_a_bits_a_mask_acc_54 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_110; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_111 = x1_a_bits_a_mask_eq_54 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_111 = x1_a_bits_a_mask_acc_54 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_111; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_112 = x1_a_bits_a_mask_eq_55 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_112 = x1_a_bits_a_mask_acc_55 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_112; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_113 = x1_a_bits_a_mask_eq_55 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_113 = x1_a_bits_a_mask_acc_55 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_113; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_114 = x1_a_bits_a_mask_eq_56 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_114 = x1_a_bits_a_mask_acc_56 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_114; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_115 = x1_a_bits_a_mask_eq_56 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_115 = x1_a_bits_a_mask_acc_56 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_115; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_116 = x1_a_bits_a_mask_eq_57 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_116 = x1_a_bits_a_mask_acc_57 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_116; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_117 = x1_a_bits_a_mask_eq_57 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_117 = x1_a_bits_a_mask_acc_57 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_117; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_118 = x1_a_bits_a_mask_eq_58 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_118 = x1_a_bits_a_mask_acc_58 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_118; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_119 = x1_a_bits_a_mask_eq_58 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_119 = x1_a_bits_a_mask_acc_58 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_119; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_120 = x1_a_bits_a_mask_eq_59 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_120 = x1_a_bits_a_mask_acc_59 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_120; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_121 = x1_a_bits_a_mask_eq_59 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_121 = x1_a_bits_a_mask_acc_59 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_121; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_122 = x1_a_bits_a_mask_eq_60 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_122 = x1_a_bits_a_mask_acc_60 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_122; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_123 = x1_a_bits_a_mask_eq_60 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_123 = x1_a_bits_a_mask_acc_60 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_123; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_124 = x1_a_bits_a_mask_eq_61 & x1_a_bits_a_mask_nbit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_124 = x1_a_bits_a_mask_acc_61 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_124; // @[Misc.scala 214:29]
  wire  x1_a_bits_a_mask_eq_125 = x1_a_bits_a_mask_eq_61 & x1_a_bits_a_mask_bit_5; // @[Misc.scala 213:27]
  wire  x1_a_bits_a_mask_acc_125 = x1_a_bits_a_mask_acc_61 | x1_a_bits_a_mask_size_5 & x1_a_bits_a_mask_eq_125; // @[Misc.scala 214:29]
  wire [7:0] x1_a_bits_a_mask_lo_lo_lo = {x1_a_bits_a_mask_acc_69,x1_a_bits_a_mask_acc_68,x1_a_bits_a_mask_acc_67,
    x1_a_bits_a_mask_acc_66,x1_a_bits_a_mask_acc_65,x1_a_bits_a_mask_acc_64,x1_a_bits_a_mask_acc_63,
    x1_a_bits_a_mask_acc_62}; // @[Cat.scala 33:92]
  wire [15:0] x1_a_bits_a_mask_lo_lo = {x1_a_bits_a_mask_acc_77,x1_a_bits_a_mask_acc_76,x1_a_bits_a_mask_acc_75,
    x1_a_bits_a_mask_acc_74,x1_a_bits_a_mask_acc_73,x1_a_bits_a_mask_acc_72,x1_a_bits_a_mask_acc_71,
    x1_a_bits_a_mask_acc_70,x1_a_bits_a_mask_lo_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] x1_a_bits_a_mask_lo_hi_lo = {x1_a_bits_a_mask_acc_85,x1_a_bits_a_mask_acc_84,x1_a_bits_a_mask_acc_83,
    x1_a_bits_a_mask_acc_82,x1_a_bits_a_mask_acc_81,x1_a_bits_a_mask_acc_80,x1_a_bits_a_mask_acc_79,
    x1_a_bits_a_mask_acc_78}; // @[Cat.scala 33:92]
  wire [31:0] x1_a_bits_a_mask_lo = {x1_a_bits_a_mask_acc_93,x1_a_bits_a_mask_acc_92,x1_a_bits_a_mask_acc_91,
    x1_a_bits_a_mask_acc_90,x1_a_bits_a_mask_acc_89,x1_a_bits_a_mask_acc_88,x1_a_bits_a_mask_acc_87,
    x1_a_bits_a_mask_acc_86,x1_a_bits_a_mask_lo_hi_lo,x1_a_bits_a_mask_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] x1_a_bits_a_mask_hi_lo_lo = {x1_a_bits_a_mask_acc_101,x1_a_bits_a_mask_acc_100,x1_a_bits_a_mask_acc_99,
    x1_a_bits_a_mask_acc_98,x1_a_bits_a_mask_acc_97,x1_a_bits_a_mask_acc_96,x1_a_bits_a_mask_acc_95,
    x1_a_bits_a_mask_acc_94}; // @[Cat.scala 33:92]
  wire [15:0] x1_a_bits_a_mask_hi_lo = {x1_a_bits_a_mask_acc_109,x1_a_bits_a_mask_acc_108,x1_a_bits_a_mask_acc_107,
    x1_a_bits_a_mask_acc_106,x1_a_bits_a_mask_acc_105,x1_a_bits_a_mask_acc_104,x1_a_bits_a_mask_acc_103,
    x1_a_bits_a_mask_acc_102,x1_a_bits_a_mask_hi_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] x1_a_bits_a_mask_hi_hi_lo = {x1_a_bits_a_mask_acc_117,x1_a_bits_a_mask_acc_116,x1_a_bits_a_mask_acc_115,
    x1_a_bits_a_mask_acc_114,x1_a_bits_a_mask_acc_113,x1_a_bits_a_mask_acc_112,x1_a_bits_a_mask_acc_111,
    x1_a_bits_a_mask_acc_110}; // @[Cat.scala 33:92]
  wire [31:0] x1_a_bits_a_mask_hi = {x1_a_bits_a_mask_acc_125,x1_a_bits_a_mask_acc_124,x1_a_bits_a_mask_acc_123,
    x1_a_bits_a_mask_acc_122,x1_a_bits_a_mask_acc_121,x1_a_bits_a_mask_acc_120,x1_a_bits_a_mask_acc_119,
    x1_a_bits_a_mask_acc_118,x1_a_bits_a_mask_hi_hi_lo,x1_a_bits_a_mask_hi_lo}; // @[Cat.scala 33:92]
  wire  _GEN_112 = 2'h1 == mem_tx_state ? reqAvailable : mem_tx_state == 2'h1; // @[CScratchpad.scala 136:19 138:24 151:23]
  wire  mem_out_a_valid = 2'h0 == mem_tx_state ? mem_tx_state == 2'h1 : _GEN_112; // @[CScratchpad.scala 136:19 138:24]
  wire  _T_13 = auto_mem_out_a_ready & mem_out_a_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_8 = 4'h0 == reqChosen ? 1'h0 : reqIdleBits_0; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_9 = 4'h1 == reqChosen ? 1'h0 : reqIdleBits_1; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_10 = 4'h2 == reqChosen ? 1'h0 : reqIdleBits_2; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_11 = 4'h3 == reqChosen ? 1'h0 : reqIdleBits_3; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_12 = 4'h4 == reqChosen ? 1'h0 : reqIdleBits_4; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_13 = 4'h5 == reqChosen ? 1'h0 : reqIdleBits_5; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_14 = 4'h6 == reqChosen ? 1'h0 : reqIdleBits_6; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_15 = 4'h7 == reqChosen ? 1'h0 : reqIdleBits_7; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_16 = 4'h8 == reqChosen ? 1'h0 : reqIdleBits_8; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_17 = 4'h9 == reqChosen ? 1'h0 : reqIdleBits_9; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_18 = 4'ha == reqChosen ? 1'h0 : reqIdleBits_10; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_19 = 4'hb == reqChosen ? 1'h0 : reqIdleBits_11; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_20 = 4'hc == reqChosen ? 1'h0 : reqIdleBits_12; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_21 = 4'hd == reqChosen ? 1'h0 : reqIdleBits_13; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_22 = 4'he == reqChosen ? 1'h0 : reqIdleBits_14; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire  _GEN_23 = 4'hf == reqChosen ? 1'h0 : reqIdleBits_15; // @[CScratchpad.scala 153:{32,32} 110:36]
  wire [33:0] _req_cache_memoryLength_T = isBelowLimit ? totalTx_memoryLength : 34'h40; // @[CScratchpad.scala 155:49]
  wire [15:0] _GEN_40 = 4'h0 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_0_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_41 = 4'h1 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_1_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_42 = 4'h2 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_2_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_43 = 4'h3 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_3_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_44 = 4'h4 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_4_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_45 = 4'h5 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_5_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_46 = 4'h6 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_6_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_47 = 4'h7 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_7_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_48 = 4'h8 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_8_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_49 = 4'h9 == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_9_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_50 = 4'ha == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_10_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_51 = 4'hb == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_11_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_52 = 4'hc == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_12_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_53 = 4'hd == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_13_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_54 = 4'he == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_14_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [15:0] _GEN_55 = 4'hf == reqChosen ? _req_cache_memoryLength_T[15:0] : req_cache_15_memoryLength; // @[CScratchpad.scala 114:30 155:{43,43}]
  wire [33:0] _totalTx_memoryLength_T_1 = totalTx_memoryLength - 34'h40; // @[CScratchpad.scala 156:54]
  wire [33:0] _totalTx_memoryAddress_T_1 = totalTx_memoryAddress + 34'h40; // @[CScratchpad.scala 158:56]
  wire [1:0] _GEN_56 = isBelowLimit ? 2'h2 : mem_tx_state; // @[CScratchpad.scala 159:28 160:24 102:37]
  wire  _GEN_57 = _T_13 ? _GEN_8 : reqIdleBits_0; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_58 = _T_13 ? _GEN_9 : reqIdleBits_1; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_59 = _T_13 ? _GEN_10 : reqIdleBits_2; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_60 = _T_13 ? _GEN_11 : reqIdleBits_3; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_61 = _T_13 ? _GEN_12 : reqIdleBits_4; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_62 = _T_13 ? _GEN_13 : reqIdleBits_5; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_63 = _T_13 ? _GEN_14 : reqIdleBits_6; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_64 = _T_13 ? _GEN_15 : reqIdleBits_7; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_65 = _T_13 ? _GEN_16 : reqIdleBits_8; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_66 = _T_13 ? _GEN_17 : reqIdleBits_9; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_67 = _T_13 ? _GEN_18 : reqIdleBits_10; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_68 = _T_13 ? _GEN_19 : reqIdleBits_11; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_69 = _T_13 ? _GEN_20 : reqIdleBits_12; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_70 = _T_13 ? _GEN_21 : reqIdleBits_13; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_71 = _T_13 ? _GEN_22 : reqIdleBits_14; // @[CScratchpad.scala 152:28 110:36]
  wire  _GEN_72 = _T_13 ? _GEN_23 : reqIdleBits_15; // @[CScratchpad.scala 152:28 110:36]
  wire [15:0] _GEN_89 = _T_13 ? _GEN_40 : req_cache_0_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_90 = _T_13 ? _GEN_41 : req_cache_1_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_91 = _T_13 ? _GEN_42 : req_cache_2_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_92 = _T_13 ? _GEN_43 : req_cache_3_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_93 = _T_13 ? _GEN_44 : req_cache_4_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_94 = _T_13 ? _GEN_45 : req_cache_5_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_95 = _T_13 ? _GEN_46 : req_cache_6_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_96 = _T_13 ? _GEN_47 : req_cache_7_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_97 = _T_13 ? _GEN_48 : req_cache_8_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_98 = _T_13 ? _GEN_49 : req_cache_9_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_99 = _T_13 ? _GEN_50 : req_cache_10_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_100 = _T_13 ? _GEN_51 : req_cache_11_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_101 = _T_13 ? _GEN_52 : req_cache_12_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_102 = _T_13 ? _GEN_53 : req_cache_13_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_103 = _T_13 ? _GEN_54 : req_cache_14_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [15:0] _GEN_104 = _T_13 ? _GEN_55 : req_cache_15_memoryLength; // @[CScratchpad.scala 152:28 114:30]
  wire [1:0] _GEN_109 = reqIdleBits_0 & reqIdleBits_1 & reqIdleBits_2 & reqIdleBits_3 & reqIdleBits_4 & reqIdleBits_5 &
    reqIdleBits_6 & reqIdleBits_7 & reqIdleBits_8 & reqIdleBits_9 & reqIdleBits_10 & reqIdleBits_11 & reqIdleBits_12 &
    reqIdleBits_13 & reqIdleBits_14 & reqIdleBits_15 ? 2'h0 : mem_tx_state; // @[CScratchpad.scala 166:40 167:22 102:37]
  wire  _GEN_113 = 2'h1 == mem_tx_state ? _GEN_57 : reqIdleBits_0; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_114 = 2'h1 == mem_tx_state ? _GEN_58 : reqIdleBits_1; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_115 = 2'h1 == mem_tx_state ? _GEN_59 : reqIdleBits_2; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_116 = 2'h1 == mem_tx_state ? _GEN_60 : reqIdleBits_3; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_117 = 2'h1 == mem_tx_state ? _GEN_61 : reqIdleBits_4; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_118 = 2'h1 == mem_tx_state ? _GEN_62 : reqIdleBits_5; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_119 = 2'h1 == mem_tx_state ? _GEN_63 : reqIdleBits_6; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_120 = 2'h1 == mem_tx_state ? _GEN_64 : reqIdleBits_7; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_121 = 2'h1 == mem_tx_state ? _GEN_65 : reqIdleBits_8; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_122 = 2'h1 == mem_tx_state ? _GEN_66 : reqIdleBits_9; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_123 = 2'h1 == mem_tx_state ? _GEN_67 : reqIdleBits_10; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_124 = 2'h1 == mem_tx_state ? _GEN_68 : reqIdleBits_11; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_125 = 2'h1 == mem_tx_state ? _GEN_69 : reqIdleBits_12; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_126 = 2'h1 == mem_tx_state ? _GEN_70 : reqIdleBits_13; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_127 = 2'h1 == mem_tx_state ? _GEN_71 : reqIdleBits_14; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_128 = 2'h1 == mem_tx_state ? _GEN_72 : reqIdleBits_15; // @[CScratchpad.scala 138:24 110:36]
  wire [15:0] _GEN_145 = 2'h1 == mem_tx_state ? _GEN_89 : req_cache_0_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_146 = 2'h1 == mem_tx_state ? _GEN_90 : req_cache_1_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_147 = 2'h1 == mem_tx_state ? _GEN_91 : req_cache_2_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_148 = 2'h1 == mem_tx_state ? _GEN_92 : req_cache_3_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_149 = 2'h1 == mem_tx_state ? _GEN_93 : req_cache_4_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_150 = 2'h1 == mem_tx_state ? _GEN_94 : req_cache_5_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_151 = 2'h1 == mem_tx_state ? _GEN_95 : req_cache_6_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_152 = 2'h1 == mem_tx_state ? _GEN_96 : req_cache_7_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_153 = 2'h1 == mem_tx_state ? _GEN_97 : req_cache_8_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_154 = 2'h1 == mem_tx_state ? _GEN_98 : req_cache_9_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_155 = 2'h1 == mem_tx_state ? _GEN_99 : req_cache_10_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_156 = 2'h1 == mem_tx_state ? _GEN_100 : req_cache_11_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_157 = 2'h1 == mem_tx_state ? _GEN_101 : req_cache_12_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_158 = 2'h1 == mem_tx_state ? _GEN_102 : req_cache_13_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_159 = 2'h1 == mem_tx_state ? _GEN_103 : req_cache_14_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_160 = 2'h1 == mem_tx_state ? _GEN_104 : req_cache_15_memoryLength; // @[CScratchpad.scala 138:24 114:30]
  wire  _GEN_171 = 2'h0 == mem_tx_state ? reqIdleBits_0 : _GEN_113; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_172 = 2'h0 == mem_tx_state ? reqIdleBits_1 : _GEN_114; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_173 = 2'h0 == mem_tx_state ? reqIdleBits_2 : _GEN_115; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_174 = 2'h0 == mem_tx_state ? reqIdleBits_3 : _GEN_116; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_175 = 2'h0 == mem_tx_state ? reqIdleBits_4 : _GEN_117; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_176 = 2'h0 == mem_tx_state ? reqIdleBits_5 : _GEN_118; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_177 = 2'h0 == mem_tx_state ? reqIdleBits_6 : _GEN_119; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_178 = 2'h0 == mem_tx_state ? reqIdleBits_7 : _GEN_120; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_179 = 2'h0 == mem_tx_state ? reqIdleBits_8 : _GEN_121; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_180 = 2'h0 == mem_tx_state ? reqIdleBits_9 : _GEN_122; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_181 = 2'h0 == mem_tx_state ? reqIdleBits_10 : _GEN_123; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_182 = 2'h0 == mem_tx_state ? reqIdleBits_11 : _GEN_124; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_183 = 2'h0 == mem_tx_state ? reqIdleBits_12 : _GEN_125; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_184 = 2'h0 == mem_tx_state ? reqIdleBits_13 : _GEN_126; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_185 = 2'h0 == mem_tx_state ? reqIdleBits_14 : _GEN_127; // @[CScratchpad.scala 138:24 110:36]
  wire  _GEN_186 = 2'h0 == mem_tx_state ? reqIdleBits_15 : _GEN_128; // @[CScratchpad.scala 138:24 110:36]
  wire [15:0] _GEN_203 = 2'h0 == mem_tx_state ? req_cache_0_memoryLength : _GEN_145; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_204 = 2'h0 == mem_tx_state ? req_cache_1_memoryLength : _GEN_146; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_205 = 2'h0 == mem_tx_state ? req_cache_2_memoryLength : _GEN_147; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_206 = 2'h0 == mem_tx_state ? req_cache_3_memoryLength : _GEN_148; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_207 = 2'h0 == mem_tx_state ? req_cache_4_memoryLength : _GEN_149; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_208 = 2'h0 == mem_tx_state ? req_cache_5_memoryLength : _GEN_150; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_209 = 2'h0 == mem_tx_state ? req_cache_6_memoryLength : _GEN_151; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_210 = 2'h0 == mem_tx_state ? req_cache_7_memoryLength : _GEN_152; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_211 = 2'h0 == mem_tx_state ? req_cache_8_memoryLength : _GEN_153; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_212 = 2'h0 == mem_tx_state ? req_cache_9_memoryLength : _GEN_154; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_213 = 2'h0 == mem_tx_state ? req_cache_10_memoryLength : _GEN_155; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_214 = 2'h0 == mem_tx_state ? req_cache_11_memoryLength : _GEN_156; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_215 = 2'h0 == mem_tx_state ? req_cache_12_memoryLength : _GEN_157; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_216 = 2'h0 == mem_tx_state ? req_cache_13_memoryLength : _GEN_158; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_217 = 2'h0 == mem_tx_state ? req_cache_14_memoryLength : _GEN_159; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_218 = 2'h0 == mem_tx_state ? req_cache_15_memoryLength : _GEN_160; // @[CScratchpad.scala 138:24 114:30]
  wire [15:0] _GEN_220 = 4'h1 == auto_mem_out_d_bits_source ? req_cache_1_memoryLength : req_cache_0_memoryLength; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_221 = 4'h2 == auto_mem_out_d_bits_source ? req_cache_2_memoryLength : _GEN_220; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_222 = 4'h3 == auto_mem_out_d_bits_source ? req_cache_3_memoryLength : _GEN_221; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_223 = 4'h4 == auto_mem_out_d_bits_source ? req_cache_4_memoryLength : _GEN_222; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_224 = 4'h5 == auto_mem_out_d_bits_source ? req_cache_5_memoryLength : _GEN_223; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_225 = 4'h6 == auto_mem_out_d_bits_source ? req_cache_6_memoryLength : _GEN_224; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_226 = 4'h7 == auto_mem_out_d_bits_source ? req_cache_7_memoryLength : _GEN_225; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_227 = 4'h8 == auto_mem_out_d_bits_source ? req_cache_8_memoryLength : _GEN_226; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_228 = 4'h9 == auto_mem_out_d_bits_source ? req_cache_9_memoryLength : _GEN_227; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_229 = 4'ha == auto_mem_out_d_bits_source ? req_cache_10_memoryLength : _GEN_228; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_230 = 4'hb == auto_mem_out_d_bits_source ? req_cache_11_memoryLength : _GEN_229; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_231 = 4'hc == auto_mem_out_d_bits_source ? req_cache_12_memoryLength : _GEN_230; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_232 = 4'hd == auto_mem_out_d_bits_source ? req_cache_13_memoryLength : _GEN_231; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_233 = 4'he == auto_mem_out_d_bits_source ? req_cache_14_memoryLength : _GEN_232; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_234 = 4'hf == auto_mem_out_d_bits_source ? req_cache_15_memoryLength : _GEN_233; // @[CScratchpad.scala 174:{40,40}]
  wire [15:0] _GEN_235 = _GEN_234 >= 16'h40 ? 16'h40 : _GEN_234; // @[CScratchpad.scala 174:55 175:39 177:39]
  wire  mem_out_d_ready = loader_io_cache_block_in_ready; // @[Nodes.scala 1212:84 CScratchpad.scala 180:19]
  wire  _T_36 = mem_out_d_ready & auto_mem_out_d_valid; // @[Decoupled.scala 51:35]
  wire [15:0] _req_cache_memoryLength_T_2 = _GEN_234 - 16'h40; // @[CScratchpad.scala 210:72]
  wire  _GEN_445 = 4'h0 == auto_mem_out_d_bits_source | _GEN_171; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_446 = 4'h1 == auto_mem_out_d_bits_source | _GEN_172; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_447 = 4'h2 == auto_mem_out_d_bits_source | _GEN_173; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_448 = 4'h3 == auto_mem_out_d_bits_source | _GEN_174; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_449 = 4'h4 == auto_mem_out_d_bits_source | _GEN_175; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_450 = 4'h5 == auto_mem_out_d_bits_source | _GEN_176; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_451 = 4'h6 == auto_mem_out_d_bits_source | _GEN_177; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_452 = 4'h7 == auto_mem_out_d_bits_source | _GEN_178; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_453 = 4'h8 == auto_mem_out_d_bits_source | _GEN_179; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_454 = 4'h9 == auto_mem_out_d_bits_source | _GEN_180; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_455 = 4'ha == auto_mem_out_d_bits_source | _GEN_181; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_456 = 4'hb == auto_mem_out_d_bits_source | _GEN_182; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_457 = 4'hc == auto_mem_out_d_bits_source | _GEN_183; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_458 = 4'hd == auto_mem_out_d_bits_source | _GEN_184; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_459 = 4'he == auto_mem_out_d_bits_source | _GEN_185; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_460 = 4'hf == auto_mem_out_d_bits_source | _GEN_186; // @[CScratchpad.scala 213:{28,28}]
  wire  _GEN_461 = _GEN_234 <= 16'h40 ? _GEN_445 : _GEN_171; // @[CScratchpad.scala 212:57]
  wire  _GEN_462 = _GEN_234 <= 16'h40 ? _GEN_446 : _GEN_172; // @[CScratchpad.scala 212:57]
  wire  _GEN_463 = _GEN_234 <= 16'h40 ? _GEN_447 : _GEN_173; // @[CScratchpad.scala 212:57]
  wire  _GEN_464 = _GEN_234 <= 16'h40 ? _GEN_448 : _GEN_174; // @[CScratchpad.scala 212:57]
  wire  _GEN_465 = _GEN_234 <= 16'h40 ? _GEN_449 : _GEN_175; // @[CScratchpad.scala 212:57]
  wire  _GEN_466 = _GEN_234 <= 16'h40 ? _GEN_450 : _GEN_176; // @[CScratchpad.scala 212:57]
  wire  _GEN_467 = _GEN_234 <= 16'h40 ? _GEN_451 : _GEN_177; // @[CScratchpad.scala 212:57]
  wire  _GEN_468 = _GEN_234 <= 16'h40 ? _GEN_452 : _GEN_178; // @[CScratchpad.scala 212:57]
  wire  _GEN_469 = _GEN_234 <= 16'h40 ? _GEN_453 : _GEN_179; // @[CScratchpad.scala 212:57]
  wire  _GEN_470 = _GEN_234 <= 16'h40 ? _GEN_454 : _GEN_180; // @[CScratchpad.scala 212:57]
  wire  _GEN_471 = _GEN_234 <= 16'h40 ? _GEN_455 : _GEN_181; // @[CScratchpad.scala 212:57]
  wire  _GEN_472 = _GEN_234 <= 16'h40 ? _GEN_456 : _GEN_182; // @[CScratchpad.scala 212:57]
  wire  _GEN_473 = _GEN_234 <= 16'h40 ? _GEN_457 : _GEN_183; // @[CScratchpad.scala 212:57]
  wire  _GEN_474 = _GEN_234 <= 16'h40 ? _GEN_458 : _GEN_184; // @[CScratchpad.scala 212:57]
  wire  _GEN_475 = _GEN_234 <= 16'h40 ? _GEN_459 : _GEN_185; // @[CScratchpad.scala 212:57]
  wire  _GEN_476 = _GEN_234 <= 16'h40 ? _GEN_460 : _GEN_186; // @[CScratchpad.scala 212:57]
  wire  _GEN_494 = _T_36 ? _GEN_461 : _GEN_171; // @[CScratchpad.scala 209:24]
  wire  _GEN_495 = _T_36 ? _GEN_462 : _GEN_172; // @[CScratchpad.scala 209:24]
  wire  _GEN_496 = _T_36 ? _GEN_463 : _GEN_173; // @[CScratchpad.scala 209:24]
  wire  _GEN_497 = _T_36 ? _GEN_464 : _GEN_174; // @[CScratchpad.scala 209:24]
  wire  _GEN_498 = _T_36 ? _GEN_465 : _GEN_175; // @[CScratchpad.scala 209:24]
  wire  _GEN_499 = _T_36 ? _GEN_466 : _GEN_176; // @[CScratchpad.scala 209:24]
  wire  _GEN_500 = _T_36 ? _GEN_467 : _GEN_177; // @[CScratchpad.scala 209:24]
  wire  _GEN_501 = _T_36 ? _GEN_468 : _GEN_178; // @[CScratchpad.scala 209:24]
  wire  _GEN_502 = _T_36 ? _GEN_469 : _GEN_179; // @[CScratchpad.scala 209:24]
  wire  _GEN_503 = _T_36 ? _GEN_470 : _GEN_180; // @[CScratchpad.scala 209:24]
  wire  _GEN_504 = _T_36 ? _GEN_471 : _GEN_181; // @[CScratchpad.scala 209:24]
  wire  _GEN_505 = _T_36 ? _GEN_472 : _GEN_182; // @[CScratchpad.scala 209:24]
  wire  _GEN_506 = _T_36 ? _GEN_473 : _GEN_183; // @[CScratchpad.scala 209:24]
  wire  _GEN_507 = _T_36 ? _GEN_474 : _GEN_184; // @[CScratchpad.scala 209:24]
  wire  _GEN_508 = _T_36 ? _GEN_475 : _GEN_185; // @[CScratchpad.scala 209:24]
  wire  _GEN_509 = _T_36 ? _GEN_476 : _GEN_186; // @[CScratchpad.scala 209:24]
  CScratchpadPackedSubwordLoader_3 loader ( // @[CScratchpad.scala 94:30]
    .clock(loader_clock),
    .reset(loader_reset),
    .io_cache_block_in_ready(loader_io_cache_block_in_ready),
    .io_cache_block_in_valid(loader_io_cache_block_in_valid),
    .io_cache_block_in_bits_len(loader_io_cache_block_in_bits_len),
    .io_sp_write_out_valid(loader_io_sp_write_out_valid)
  );
  assign auto_mem_out_a_valid = 2'h0 == mem_tx_state ? mem_tx_state == 2'h1 : _GEN_112; // @[CScratchpad.scala 136:19 138:24]
  assign auto_mem_out_a_bits_size = txEmitLengthLg[2:0]; // @[Edges.scala 447:17 450:15]
  assign auto_mem_out_a_bits_source = reqIdleBits_0 ? 4'h0 : _reqChosen_T_13; // @[Mux.scala 47:70]
  assign auto_mem_out_a_bits_address = totalTx_memoryAddress; // @[Edges.scala 447:17 452:15]
  assign auto_mem_out_a_bits_mask = {x1_a_bits_a_mask_hi,x1_a_bits_a_mask_lo}; // @[Cat.scala 33:92]
  assign auto_mem_out_d_ready = loader_io_cache_block_in_ready; // @[Nodes.scala 1212:84 CScratchpad.scala 180:19]
  assign loader_clock = clock;
  assign loader_reset = reset;
  assign loader_io_cache_block_in_valid = auto_mem_out_d_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign loader_io_cache_block_in_bits_len = _GEN_235[6:0];
  always @(posedge clock) begin
    if (reset) begin // @[CScratchpad.scala 102:37]
      mem_tx_state <= 2'h0; // @[CScratchpad.scala 102:37]
    end else if (!(2'h0 == mem_tx_state)) begin // @[CScratchpad.scala 138:24]
      if (2'h1 == mem_tx_state) begin // @[CScratchpad.scala 138:24]
        if (_T_13) begin // @[CScratchpad.scala 152:28]
          mem_tx_state <= _GEN_56;
        end
      end else if (2'h2 == mem_tx_state) begin // @[CScratchpad.scala 138:24]
        mem_tx_state <= _GEN_109;
      end
    end
    reqIdleBits_0 <= reset | _GEN_494; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_1 <= reset | _GEN_495; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_2 <= reset | _GEN_496; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_3 <= reset | _GEN_497; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_4 <= reset | _GEN_498; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_5 <= reset | _GEN_499; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_6 <= reset | _GEN_500; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_7 <= reset | _GEN_501; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_8 <= reset | _GEN_502; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_9 <= reset | _GEN_503; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_10 <= reset | _GEN_504; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_11 <= reset | _GEN_505; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_12 <= reset | _GEN_506; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_13 <= reset | _GEN_507; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_14 <= reset | _GEN_508; // @[CScratchpad.scala 110:{36,36}]
    reqIdleBits_15 <= reset | _GEN_509; // @[CScratchpad.scala 110:{36,36}]
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h0 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_0_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_0_memoryLength <= _GEN_203;
      end
    end else begin
      req_cache_0_memoryLength <= _GEN_203;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h1 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_1_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_1_memoryLength <= _GEN_204;
      end
    end else begin
      req_cache_1_memoryLength <= _GEN_204;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h2 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_2_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_2_memoryLength <= _GEN_205;
      end
    end else begin
      req_cache_2_memoryLength <= _GEN_205;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h3 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_3_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_3_memoryLength <= _GEN_206;
      end
    end else begin
      req_cache_3_memoryLength <= _GEN_206;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h4 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_4_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_4_memoryLength <= _GEN_207;
      end
    end else begin
      req_cache_4_memoryLength <= _GEN_207;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h5 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_5_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_5_memoryLength <= _GEN_208;
      end
    end else begin
      req_cache_5_memoryLength <= _GEN_208;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h6 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_6_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_6_memoryLength <= _GEN_209;
      end
    end else begin
      req_cache_6_memoryLength <= _GEN_209;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h7 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_7_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_7_memoryLength <= _GEN_210;
      end
    end else begin
      req_cache_7_memoryLength <= _GEN_210;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h8 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_8_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_8_memoryLength <= _GEN_211;
      end
    end else begin
      req_cache_8_memoryLength <= _GEN_211;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'h9 == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_9_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_9_memoryLength <= _GEN_212;
      end
    end else begin
      req_cache_9_memoryLength <= _GEN_212;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'ha == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_10_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_10_memoryLength <= _GEN_213;
      end
    end else begin
      req_cache_10_memoryLength <= _GEN_213;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'hb == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_11_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_11_memoryLength <= _GEN_214;
      end
    end else begin
      req_cache_11_memoryLength <= _GEN_214;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'hc == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_12_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_12_memoryLength <= _GEN_215;
      end
    end else begin
      req_cache_12_memoryLength <= _GEN_215;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'hd == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_13_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_13_memoryLength <= _GEN_216;
      end
    end else begin
      req_cache_13_memoryLength <= _GEN_216;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'he == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_14_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_14_memoryLength <= _GEN_217;
      end
    end else begin
      req_cache_14_memoryLength <= _GEN_217;
    end
    if (_T_36) begin // @[CScratchpad.scala 209:24]
      if (4'hf == auto_mem_out_d_bits_source) begin // @[CScratchpad.scala 210:37]
        req_cache_15_memoryLength <= _req_cache_memoryLength_T_2; // @[CScratchpad.scala 210:37]
      end else begin
        req_cache_15_memoryLength <= _GEN_218;
      end
    end else begin
      req_cache_15_memoryLength <= _GEN_218;
    end
    if (!(2'h0 == mem_tx_state)) begin // @[CScratchpad.scala 138:24]
      if (2'h1 == mem_tx_state) begin // @[CScratchpad.scala 138:24]
        if (_T_13) begin // @[CScratchpad.scala 152:28]
          totalTx_memoryAddress <= _totalTx_memoryAddress_T_1; // @[CScratchpad.scala 158:31]
        end
      end
    end
    if (!(2'h0 == mem_tx_state)) begin // @[CScratchpad.scala 138:24]
      if (2'h1 == mem_tx_state) begin // @[CScratchpad.scala 138:24]
        if (_T_13) begin // @[CScratchpad.scala 152:28]
          totalTx_memoryLength <= _totalTx_memoryLength_T_1; // @[CScratchpad.scala 156:30]
        end
      end
    end
  end
endmodule
module SequentialWriter(
  input          clock,
  input          reset,
  output         io_req_ready,
  input          io_req_valid,
  input  [33:0]  io_req_bits_addr,
  input  [33:0]  io_req_bits_len,
  output         io_channel_data_ready,
  input          io_channel_data_valid,
  input  [31:0]  io_channel_data_bits,
  output         io_channel_channelIdle,
  input          tl_out_a_ready,
  output         tl_out_a_valid,
  output         tl_out_a_bits_source,
  output [33:0]  tl_out_a_bits_address,
  output [63:0]  tl_out_a_bits_mask,
  output [511:0] tl_out_a_bits_data,
  output         tl_out_d_ready,
  input          tl_out_d_valid,
  input          tl_out_d_bits_source
);
  reg [1:0] state; // @[Writers.scala 36:30]
  reg  txStates_0; // @[Writers.scala 42:33]
  reg  txStates_1; // @[Writers.scala 42:33]
  wire  _txPriority_T = ~txStates_0; // @[Writers.scala 43:62]
  wire  _txPriority_T_1 = ~txStates_1; // @[Writers.scala 43:62]
  wire [1:0] _txPriority_enc_T = _txPriority_T_1 ? 2'h2 : 2'h0; // @[Mux.scala 47:70]
  wire [1:0] txPriority_enc = _txPriority_T ? 2'h1 : _txPriority_enc_T; // @[Mux.scala 47:70]
  wire  txPriority_0 = txPriority_enc[0]; // @[OneHot.scala 82:30]
  wire  txPriority_1 = txPriority_enc[1]; // @[OneHot.scala 82:30]
  wire  haveTransactionToDo = txStates_0 | txStates_1; // @[Writers.scala 45:80]
  wire  haveAvailableTxSlot = _txPriority_T | _txPriority_T_1; // @[Writers.scala 46:78]
  reg [27:0] addr; // @[Writers.scala 57:25]
  reg [31:0] req_len; // @[Writers.scala 60:28]
  wire [27:0] nextAddr = addr + 28'h1; // @[Writers.scala 64:31]
  reg [3:0] idx; // @[Writers.scala 66:24]
  reg [31:0] dataBuf_0; // @[Writers.scala 68:28]
  reg [31:0] dataBuf_1; // @[Writers.scala 68:28]
  reg [31:0] dataBuf_2; // @[Writers.scala 68:28]
  reg [31:0] dataBuf_3; // @[Writers.scala 68:28]
  reg [31:0] dataBuf_4; // @[Writers.scala 68:28]
  reg [31:0] dataBuf_5; // @[Writers.scala 68:28]
  reg [31:0] dataBuf_6; // @[Writers.scala 68:28]
  reg [31:0] dataBuf_7; // @[Writers.scala 68:28]
  reg [31:0] dataBuf_8; // @[Writers.scala 68:28]
  reg [31:0] dataBuf_9; // @[Writers.scala 68:28]
  reg [31:0] dataBuf_10; // @[Writers.scala 68:28]
  reg [31:0] dataBuf_11; // @[Writers.scala 68:28]
  reg [31:0] dataBuf_12; // @[Writers.scala 68:28]
  reg [31:0] dataBuf_13; // @[Writers.scala 68:28]
  reg [31:0] dataBuf_14; // @[Writers.scala 68:28]
  reg [31:0] dataBuf_15; // @[Writers.scala 68:28]
  reg [15:0] dataValid; // @[Writers.scala 69:30]
  wire [255:0] wdata_lo = {dataBuf_7,dataBuf_6,dataBuf_5,dataBuf_4,dataBuf_3,dataBuf_2,dataBuf_1,dataBuf_0}; // @[Writers.scala 71:31]
  wire [255:0] wdata_hi = {dataBuf_15,dataBuf_14,dataBuf_13,dataBuf_12,dataBuf_11,dataBuf_10,dataBuf_9,dataBuf_8}; // @[Writers.scala 71:31]
  wire [3:0] _wmask_T_17 = dataValid[0] ? 4'hf : 4'h0; // @[Bitwise.scala 77:12]
  wire [3:0] _wmask_T_19 = dataValid[1] ? 4'hf : 4'h0; // @[Bitwise.scala 77:12]
  wire [3:0] _wmask_T_21 = dataValid[2] ? 4'hf : 4'h0; // @[Bitwise.scala 77:12]
  wire [3:0] _wmask_T_23 = dataValid[3] ? 4'hf : 4'h0; // @[Bitwise.scala 77:12]
  wire [3:0] _wmask_T_25 = dataValid[4] ? 4'hf : 4'h0; // @[Bitwise.scala 77:12]
  wire [3:0] _wmask_T_27 = dataValid[5] ? 4'hf : 4'h0; // @[Bitwise.scala 77:12]
  wire [3:0] _wmask_T_29 = dataValid[6] ? 4'hf : 4'h0; // @[Bitwise.scala 77:12]
  wire [3:0] _wmask_T_31 = dataValid[7] ? 4'hf : 4'h0; // @[Bitwise.scala 77:12]
  wire [3:0] _wmask_T_33 = dataValid[8] ? 4'hf : 4'h0; // @[Bitwise.scala 77:12]
  wire [3:0] _wmask_T_35 = dataValid[9] ? 4'hf : 4'h0; // @[Bitwise.scala 77:12]
  wire [3:0] _wmask_T_37 = dataValid[10] ? 4'hf : 4'h0; // @[Bitwise.scala 77:12]
  wire [3:0] _wmask_T_39 = dataValid[11] ? 4'hf : 4'h0; // @[Bitwise.scala 77:12]
  wire [3:0] _wmask_T_41 = dataValid[12] ? 4'hf : 4'h0; // @[Bitwise.scala 77:12]
  wire [3:0] _wmask_T_43 = dataValid[13] ? 4'hf : 4'h0; // @[Bitwise.scala 77:12]
  wire [3:0] _wmask_T_45 = dataValid[14] ? 4'hf : 4'h0; // @[Bitwise.scala 77:12]
  wire [3:0] _wmask_T_47 = dataValid[15] ? 4'hf : 4'h0; // @[Bitwise.scala 77:12]
  wire [31:0] wmask_lo = {_wmask_T_31,_wmask_T_29,_wmask_T_27,_wmask_T_25,_wmask_T_23,_wmask_T_21,_wmask_T_19,
    _wmask_T_17}; // @[Cat.scala 33:92]
  wire [31:0] wmask_hi = {_wmask_T_47,_wmask_T_45,_wmask_T_43,_wmask_T_41,_wmask_T_39,_wmask_T_37,_wmask_T_35,
    _wmask_T_33}; // @[Cat.scala 33:92]
  reg  allocatedTransaction; // @[Writers.scala 74:45]
  wire  _T = tl_out_d_ready & tl_out_d_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_0 = ~tl_out_d_bits_source ? 1'h0 : txStates_0; // @[Writers.scala 42:33 82:{36,36}]
  wire  _GEN_1 = tl_out_d_bits_source ? 1'h0 : txStates_1; // @[Writers.scala 42:33 82:{36,36}]
  wire  _GEN_2 = _T ? _GEN_0 : txStates_0; // @[Writers.scala 81:23 42:33]
  wire  _GEN_3 = _T ? _GEN_1 : txStates_1; // @[Writers.scala 81:23 42:33]
  wire  _T_1 = 2'h0 == state; // @[Writers.scala 85:17]
  wire  _T_2 = io_req_ready & io_req_valid; // @[Decoupled.scala 51:35]
  wire [4:0] _GEN_4 = _T_2 ? io_req_bits_addr[6:2] : {{1'd0}, idx}; // @[Writers.scala 87:25 91:15 66:24]
  wire  _T_9 = io_channel_data_ready & io_channel_data_valid; // @[Decoupled.scala 51:35]
  wire [15:0] _dataValid_T = 16'h1 << idx; // @[OneHot.scala 57:35]
  wire [15:0] _dataValid_T_1 = dataValid | _dataValid_T; // @[Writers.scala 110:32]
  wire [3:0] _idx_T_2 = idx + 4'h1; // @[Writers.scala 111:20]
  wire [31:0] _req_len_T_2 = req_len - 32'h1; // @[Writers.scala 112:28]
  wire [1:0] _GEN_25 = idx == 4'hf | req_len == 32'h1 ? 2'h2 : state; // @[Writers.scala 113:63 114:17 36:30]
  wire [3:0] _GEN_43 = _T_9 ? _idx_T_2 : idx; // @[Writers.scala 108:34 111:13 66:24]
  wire [1:0] _allocatedTransaction_T = {txPriority_1,txPriority_0}; // @[Cat.scala 33:92]
  wire  _GEN_46 = haveAvailableTxSlot ? _allocatedTransaction_T[1] : allocatedTransaction; // @[Writers.scala 119:33 120:30 74:45]
  wire [1:0] _GEN_47 = haveAvailableTxSlot ? 2'h3 : state; // @[Writers.scala 119:33 121:15 36:30]
  wire  _T_15 = tl_out_a_ready & tl_out_a_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_48 = ~allocatedTransaction | _GEN_2; // @[Writers.scala 135:{40,40}]
  wire  _GEN_49 = allocatedTransaction | _GEN_3; // @[Writers.scala 135:{40,40}]
  wire [1:0] _GEN_50 = req_len == 32'h0 ? 2'h0 : 2'h1; // @[Writers.scala 139:46 140:17 143:17]
  wire  _GEN_52 = _T_15 ? _GEN_48 : _GEN_2; // @[Writers.scala 134:27]
  wire  _GEN_53 = _T_15 ? _GEN_49 : _GEN_3; // @[Writers.scala 134:27]
  wire [27:0] _GEN_54 = _T_15 ? nextAddr : addr; // @[Writers.scala 134:27 136:14 57:25]
  wire [3:0] _GEN_55 = _T_15 ? 4'h0 : idx; // @[Writers.scala 134:27 137:13 66:24]
  wire [15:0] _GEN_56 = _T_15 ? 16'h0 : dataValid; // @[Writers.scala 134:27 138:19 69:30]
  wire [1:0] _GEN_57 = _T_15 ? _GEN_50 : state; // @[Writers.scala 134:27 36:30]
  wire  _GEN_68 = 2'h3 == state ? _GEN_52 : _GEN_2; // @[Writers.scala 85:17]
  wire  _GEN_69 = 2'h3 == state ? _GEN_53 : _GEN_3; // @[Writers.scala 85:17]
  wire [3:0] _GEN_71 = 2'h3 == state ? _GEN_55 : idx; // @[Writers.scala 85:17 66:24]
  wire [1:0] _GEN_73 = 2'h3 == state ? _GEN_57 : state; // @[Writers.scala 85:17 36:30]
  wire  _GEN_77 = 2'h2 == state ? 1'h0 : 2'h3 == state; // @[Writers.scala 85:17 78:18]
  wire [3:0] _GEN_89 = 2'h2 == state ? idx : _GEN_71; // @[Writers.scala 85:17 66:24]
  wire [3:0] _GEN_109 = 2'h1 == state ? _GEN_43 : _GEN_89; // @[Writers.scala 85:17]
  wire  _GEN_113 = 2'h1 == state ? 1'h0 : _GEN_77; // @[Writers.scala 85:17 78:18]
  wire [4:0] _GEN_126 = 2'h0 == state ? _GEN_4 : {{1'd0}, _GEN_109}; // @[Writers.scala 85:17]
  assign io_req_ready = state == 2'h0; // @[Writers.scala 149:25]
  assign io_channel_data_ready = state == 2'h1; // @[Writers.scala 150:34]
  assign io_channel_channelIdle = ~haveTransactionToDo; // @[Writers.scala 49:29]
  assign tl_out_a_valid = 2'h0 == state ? 1'h0 : _GEN_113; // @[Writers.scala 85:17 78:18]
  assign tl_out_a_bits_source = allocatedTransaction; // @[Edges.scala 483:17 487:15]
  assign tl_out_a_bits_address = {addr,6'h0}; // @[Cat.scala 33:92]
  assign tl_out_a_bits_mask = {wmask_hi,wmask_lo}; // @[Cat.scala 33:92]
  assign tl_out_a_bits_data = {wdata_hi,wdata_lo}; // @[Writers.scala 71:31]
  assign tl_out_d_ready = txStates_0 | txStates_1; // @[Writers.scala 45:80]
  always @(posedge clock) begin
    if (reset) begin // @[Writers.scala 36:30]
      state <= 2'h0; // @[Writers.scala 36:30]
    end else if (2'h0 == state) begin // @[Writers.scala 85:17]
      if (_T_2) begin // @[Writers.scala 87:25]
        state <= 2'h1; // @[Writers.scala 102:15]
      end
    end else if (2'h1 == state) begin // @[Writers.scala 85:17]
      if (_T_9) begin // @[Writers.scala 108:34]
        state <= _GEN_25;
      end
    end else if (2'h2 == state) begin // @[Writers.scala 85:17]
      state <= _GEN_47;
    end else begin
      state <= _GEN_73;
    end
    if (reset) begin // @[Writers.scala 42:33]
      txStates_0 <= 1'h0; // @[Writers.scala 42:33]
    end else if (2'h0 == state) begin // @[Writers.scala 85:17]
      txStates_0 <= _GEN_2;
    end else if (2'h1 == state) begin // @[Writers.scala 85:17]
      txStates_0 <= _GEN_2;
    end else if (2'h2 == state) begin // @[Writers.scala 85:17]
      txStates_0 <= _GEN_2;
    end else begin
      txStates_0 <= _GEN_68;
    end
    if (reset) begin // @[Writers.scala 42:33]
      txStates_1 <= 1'h0; // @[Writers.scala 42:33]
    end else if (2'h0 == state) begin // @[Writers.scala 85:17]
      txStates_1 <= _GEN_3;
    end else if (2'h1 == state) begin // @[Writers.scala 85:17]
      txStates_1 <= _GEN_3;
    end else if (2'h2 == state) begin // @[Writers.scala 85:17]
      txStates_1 <= _GEN_3;
    end else begin
      txStates_1 <= _GEN_69;
    end
    if (2'h0 == state) begin // @[Writers.scala 85:17]
      if (_T_2) begin // @[Writers.scala 87:25]
        addr <= io_req_bits_addr[33:6]; // @[Writers.scala 94:14]
      end
    end else if (!(2'h1 == state)) begin // @[Writers.scala 85:17]
      if (!(2'h2 == state)) begin // @[Writers.scala 85:17]
        if (2'h3 == state) begin // @[Writers.scala 85:17]
          addr <= _GEN_54;
        end
      end
    end
    if (2'h0 == state) begin // @[Writers.scala 85:17]
      if (_T_2) begin // @[Writers.scala 87:25]
        req_len <= io_req_bits_len[33:2]; // @[Writers.scala 93:17]
      end
    end else if (2'h1 == state) begin // @[Writers.scala 85:17]
      if (_T_9) begin // @[Writers.scala 108:34]
        req_len <= _req_len_T_2; // @[Writers.scala 112:17]
      end
    end
    idx <= _GEN_126[3:0];
    if (!(2'h0 == state)) begin // @[Writers.scala 85:17]
      if (2'h1 == state) begin // @[Writers.scala 85:17]
        if (_T_9) begin // @[Writers.scala 108:34]
          if (4'h0 == idx) begin // @[Writers.scala 109:22]
            dataBuf_0 <= io_channel_data_bits; // @[Writers.scala 109:22]
          end
        end
      end
    end
    if (!(2'h0 == state)) begin // @[Writers.scala 85:17]
      if (2'h1 == state) begin // @[Writers.scala 85:17]
        if (_T_9) begin // @[Writers.scala 108:34]
          if (4'h1 == idx) begin // @[Writers.scala 109:22]
            dataBuf_1 <= io_channel_data_bits; // @[Writers.scala 109:22]
          end
        end
      end
    end
    if (!(2'h0 == state)) begin // @[Writers.scala 85:17]
      if (2'h1 == state) begin // @[Writers.scala 85:17]
        if (_T_9) begin // @[Writers.scala 108:34]
          if (4'h2 == idx) begin // @[Writers.scala 109:22]
            dataBuf_2 <= io_channel_data_bits; // @[Writers.scala 109:22]
          end
        end
      end
    end
    if (!(2'h0 == state)) begin // @[Writers.scala 85:17]
      if (2'h1 == state) begin // @[Writers.scala 85:17]
        if (_T_9) begin // @[Writers.scala 108:34]
          if (4'h3 == idx) begin // @[Writers.scala 109:22]
            dataBuf_3 <= io_channel_data_bits; // @[Writers.scala 109:22]
          end
        end
      end
    end
    if (!(2'h0 == state)) begin // @[Writers.scala 85:17]
      if (2'h1 == state) begin // @[Writers.scala 85:17]
        if (_T_9) begin // @[Writers.scala 108:34]
          if (4'h4 == idx) begin // @[Writers.scala 109:22]
            dataBuf_4 <= io_channel_data_bits; // @[Writers.scala 109:22]
          end
        end
      end
    end
    if (!(2'h0 == state)) begin // @[Writers.scala 85:17]
      if (2'h1 == state) begin // @[Writers.scala 85:17]
        if (_T_9) begin // @[Writers.scala 108:34]
          if (4'h5 == idx) begin // @[Writers.scala 109:22]
            dataBuf_5 <= io_channel_data_bits; // @[Writers.scala 109:22]
          end
        end
      end
    end
    if (!(2'h0 == state)) begin // @[Writers.scala 85:17]
      if (2'h1 == state) begin // @[Writers.scala 85:17]
        if (_T_9) begin // @[Writers.scala 108:34]
          if (4'h6 == idx) begin // @[Writers.scala 109:22]
            dataBuf_6 <= io_channel_data_bits; // @[Writers.scala 109:22]
          end
        end
      end
    end
    if (!(2'h0 == state)) begin // @[Writers.scala 85:17]
      if (2'h1 == state) begin // @[Writers.scala 85:17]
        if (_T_9) begin // @[Writers.scala 108:34]
          if (4'h7 == idx) begin // @[Writers.scala 109:22]
            dataBuf_7 <= io_channel_data_bits; // @[Writers.scala 109:22]
          end
        end
      end
    end
    if (!(2'h0 == state)) begin // @[Writers.scala 85:17]
      if (2'h1 == state) begin // @[Writers.scala 85:17]
        if (_T_9) begin // @[Writers.scala 108:34]
          if (4'h8 == idx) begin // @[Writers.scala 109:22]
            dataBuf_8 <= io_channel_data_bits; // @[Writers.scala 109:22]
          end
        end
      end
    end
    if (!(2'h0 == state)) begin // @[Writers.scala 85:17]
      if (2'h1 == state) begin // @[Writers.scala 85:17]
        if (_T_9) begin // @[Writers.scala 108:34]
          if (4'h9 == idx) begin // @[Writers.scala 109:22]
            dataBuf_9 <= io_channel_data_bits; // @[Writers.scala 109:22]
          end
        end
      end
    end
    if (!(2'h0 == state)) begin // @[Writers.scala 85:17]
      if (2'h1 == state) begin // @[Writers.scala 85:17]
        if (_T_9) begin // @[Writers.scala 108:34]
          if (4'ha == idx) begin // @[Writers.scala 109:22]
            dataBuf_10 <= io_channel_data_bits; // @[Writers.scala 109:22]
          end
        end
      end
    end
    if (!(2'h0 == state)) begin // @[Writers.scala 85:17]
      if (2'h1 == state) begin // @[Writers.scala 85:17]
        if (_T_9) begin // @[Writers.scala 108:34]
          if (4'hb == idx) begin // @[Writers.scala 109:22]
            dataBuf_11 <= io_channel_data_bits; // @[Writers.scala 109:22]
          end
        end
      end
    end
    if (!(2'h0 == state)) begin // @[Writers.scala 85:17]
      if (2'h1 == state) begin // @[Writers.scala 85:17]
        if (_T_9) begin // @[Writers.scala 108:34]
          if (4'hc == idx) begin // @[Writers.scala 109:22]
            dataBuf_12 <= io_channel_data_bits; // @[Writers.scala 109:22]
          end
        end
      end
    end
    if (!(2'h0 == state)) begin // @[Writers.scala 85:17]
      if (2'h1 == state) begin // @[Writers.scala 85:17]
        if (_T_9) begin // @[Writers.scala 108:34]
          if (4'hd == idx) begin // @[Writers.scala 109:22]
            dataBuf_13 <= io_channel_data_bits; // @[Writers.scala 109:22]
          end
        end
      end
    end
    if (!(2'h0 == state)) begin // @[Writers.scala 85:17]
      if (2'h1 == state) begin // @[Writers.scala 85:17]
        if (_T_9) begin // @[Writers.scala 108:34]
          if (4'he == idx) begin // @[Writers.scala 109:22]
            dataBuf_14 <= io_channel_data_bits; // @[Writers.scala 109:22]
          end
        end
      end
    end
    if (!(2'h0 == state)) begin // @[Writers.scala 85:17]
      if (2'h1 == state) begin // @[Writers.scala 85:17]
        if (_T_9) begin // @[Writers.scala 108:34]
          if (4'hf == idx) begin // @[Writers.scala 109:22]
            dataBuf_15 <= io_channel_data_bits; // @[Writers.scala 109:22]
          end
        end
      end
    end
    if (2'h0 == state) begin // @[Writers.scala 85:17]
      if (_T_2) begin // @[Writers.scala 87:25]
        dataValid <= 16'h0; // @[Writers.scala 95:19]
      end
    end else if (2'h1 == state) begin // @[Writers.scala 85:17]
      if (_T_9) begin // @[Writers.scala 108:34]
        dataValid <= _dataValid_T_1; // @[Writers.scala 110:19]
      end
    end else if (!(2'h2 == state)) begin // @[Writers.scala 85:17]
      if (2'h3 == state) begin // @[Writers.scala 85:17]
        dataValid <= _GEN_56;
      end
    end
    if (reset) begin // @[Writers.scala 74:45]
      allocatedTransaction <= 1'h0; // @[Writers.scala 74:45]
    end else if (!(2'h0 == state)) begin // @[Writers.scala 85:17]
      if (!(2'h1 == state)) begin // @[Writers.scala 85:17]
        if (2'h2 == state) begin // @[Writers.scala 85:17]
          allocatedTransaction <= _GEN_46;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1 & _T_2 & ~reset & ~(io_req_bits_addr[1:0] == 2'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed: FixedSequentialWriteChannel: Unaligned request\n    at Writers.scala:98 assert(io.req.bits.addr(log2Ceil(nBytes) - 1, 0) === 0.U,\n"
            ); // @[Writers.scala 98:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(io_req_bits_addr[1:0] == 2'h0) & (_T_1 & _T_2 & ~reset)) begin
          $fatal; // @[Writers.scala 98:17]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComposerCoreWrapper(
  input          clock,
  input          reset,
  input          auto_solvated_mem_out_a_ready,
  output         auto_solvated_mem_out_a_valid,
  output [2:0]   auto_solvated_mem_out_a_bits_size,
  output [3:0]   auto_solvated_mem_out_a_bits_source,
  output [33:0]  auto_solvated_mem_out_a_bits_address,
  output [63:0]  auto_solvated_mem_out_a_bits_mask,
  output         auto_solvated_mem_out_d_ready,
  input          auto_solvated_mem_out_d_valid,
  input  [3:0]   auto_solvated_mem_out_d_bits_source,
  input          auto_nonBonded_mem_out_a_ready,
  output         auto_nonBonded_mem_out_a_valid,
  output [2:0]   auto_nonBonded_mem_out_a_bits_size,
  output [3:0]   auto_nonBonded_mem_out_a_bits_source,
  output [33:0]  auto_nonBonded_mem_out_a_bits_address,
  output [63:0]  auto_nonBonded_mem_out_a_bits_mask,
  output         auto_nonBonded_mem_out_d_ready,
  input          auto_nonBonded_mem_out_d_valid,
  input  [3:0]   auto_nonBonded_mem_out_d_bits_source,
  input          auto_halfNonBonded_mem_out_a_ready,
  output         auto_halfNonBonded_mem_out_a_valid,
  output [2:0]   auto_halfNonBonded_mem_out_a_bits_size,
  output [3:0]   auto_halfNonBonded_mem_out_a_bits_source,
  output [33:0]  auto_halfNonBonded_mem_out_a_bits_address,
  output [63:0]  auto_halfNonBonded_mem_out_a_bits_mask,
  output         auto_halfNonBonded_mem_out_d_ready,
  input          auto_halfNonBonded_mem_out_d_valid,
  input  [3:0]   auto_halfNonBonded_mem_out_d_bits_source,
  input          auto_data_mem_out_a_ready,
  output         auto_data_mem_out_a_valid,
  output [2:0]   auto_data_mem_out_a_bits_size,
  output [3:0]   auto_data_mem_out_a_bits_source,
  output [33:0]  auto_data_mem_out_a_bits_address,
  output [63:0]  auto_data_mem_out_a_bits_mask,
  output         auto_data_mem_out_d_ready,
  input          auto_data_mem_out_d_valid,
  input  [3:0]   auto_data_mem_out_d_bits_source,
  input  [511:0] auto_data_mem_out_d_bits_data,
  input          auto_writers_out_a_ready,
  output         auto_writers_out_a_valid,
  output         auto_writers_out_a_bits_source,
  output [33:0]  auto_writers_out_a_bits_address,
  output [63:0]  auto_writers_out_a_bits_mask,
  output [511:0] auto_writers_out_a_bits_data,
  output         auto_writers_out_d_ready,
  input          auto_writers_out_d_valid,
  input          auto_writers_out_d_bits_source,
  output         io_req_ready,
  input          io_req_valid,
  input  [4:0]   io_req_bits_inst_rs1,
  input  [55:0]  io_req_bits_payload1,
  input  [63:0]  io_req_bits_payload2,
  input          io_resp_ready,
  output         io_resp_valid,
  input          myWriters_WriteChannel_valid,
  input  [33:0]  myWriters_WriteChannel_bits_addr,
  input  [33:0]  myWriters_WriteChannel_bits_len
);
  wire  data_clock; // @[ComposerCore.scala 76:32]
  wire  data_reset; // @[ComposerCore.scala 76:32]
  wire  data_auto_mem_out_a_ready; // @[ComposerCore.scala 76:32]
  wire  data_auto_mem_out_a_valid; // @[ComposerCore.scala 76:32]
  wire [2:0] data_auto_mem_out_a_bits_size; // @[ComposerCore.scala 76:32]
  wire [3:0] data_auto_mem_out_a_bits_source; // @[ComposerCore.scala 76:32]
  wire [33:0] data_auto_mem_out_a_bits_address; // @[ComposerCore.scala 76:32]
  wire [63:0] data_auto_mem_out_a_bits_mask; // @[ComposerCore.scala 76:32]
  wire  data_auto_mem_out_d_ready; // @[ComposerCore.scala 76:32]
  wire  data_auto_mem_out_d_valid; // @[ComposerCore.scala 76:32]
  wire [3:0] data_auto_mem_out_d_bits_source; // @[ComposerCore.scala 76:32]
  wire [511:0] data_auto_mem_out_d_bits_data; // @[ComposerCore.scala 76:32]
  wire  data_access_readReq_valid; // @[ComposerCore.scala 76:32]
  wire  data_access_readRes_valid; // @[ComposerCore.scala 76:32]
  wire [127:0] data_access_readRes_bits; // @[ComposerCore.scala 76:32]
  wire  halfNonBonded_clock; // @[ComposerCore.scala 76:32]
  wire  halfNonBonded_reset; // @[ComposerCore.scala 76:32]
  wire  halfNonBonded_auto_mem_out_a_ready; // @[ComposerCore.scala 76:32]
  wire  halfNonBonded_auto_mem_out_a_valid; // @[ComposerCore.scala 76:32]
  wire [2:0] halfNonBonded_auto_mem_out_a_bits_size; // @[ComposerCore.scala 76:32]
  wire [3:0] halfNonBonded_auto_mem_out_a_bits_source; // @[ComposerCore.scala 76:32]
  wire [33:0] halfNonBonded_auto_mem_out_a_bits_address; // @[ComposerCore.scala 76:32]
  wire [63:0] halfNonBonded_auto_mem_out_a_bits_mask; // @[ComposerCore.scala 76:32]
  wire  halfNonBonded_auto_mem_out_d_ready; // @[ComposerCore.scala 76:32]
  wire  halfNonBonded_auto_mem_out_d_valid; // @[ComposerCore.scala 76:32]
  wire [3:0] halfNonBonded_auto_mem_out_d_bits_source; // @[ComposerCore.scala 76:32]
  wire  nonBonded_clock; // @[ComposerCore.scala 76:32]
  wire  nonBonded_reset; // @[ComposerCore.scala 76:32]
  wire  nonBonded_auto_mem_out_a_ready; // @[ComposerCore.scala 76:32]
  wire  nonBonded_auto_mem_out_a_valid; // @[ComposerCore.scala 76:32]
  wire [2:0] nonBonded_auto_mem_out_a_bits_size; // @[ComposerCore.scala 76:32]
  wire [3:0] nonBonded_auto_mem_out_a_bits_source; // @[ComposerCore.scala 76:32]
  wire [33:0] nonBonded_auto_mem_out_a_bits_address; // @[ComposerCore.scala 76:32]
  wire [63:0] nonBonded_auto_mem_out_a_bits_mask; // @[ComposerCore.scala 76:32]
  wire  nonBonded_auto_mem_out_d_ready; // @[ComposerCore.scala 76:32]
  wire  nonBonded_auto_mem_out_d_valid; // @[ComposerCore.scala 76:32]
  wire [3:0] nonBonded_auto_mem_out_d_bits_source; // @[ComposerCore.scala 76:32]
  wire  solvated_clock; // @[ComposerCore.scala 76:32]
  wire  solvated_reset; // @[ComposerCore.scala 76:32]
  wire  solvated_auto_mem_out_a_ready; // @[ComposerCore.scala 76:32]
  wire  solvated_auto_mem_out_a_valid; // @[ComposerCore.scala 76:32]
  wire [2:0] solvated_auto_mem_out_a_bits_size; // @[ComposerCore.scala 76:32]
  wire [3:0] solvated_auto_mem_out_a_bits_source; // @[ComposerCore.scala 76:32]
  wire [33:0] solvated_auto_mem_out_a_bits_address; // @[ComposerCore.scala 76:32]
  wire [63:0] solvated_auto_mem_out_a_bits_mask; // @[ComposerCore.scala 76:32]
  wire  solvated_auto_mem_out_d_ready; // @[ComposerCore.scala 76:32]
  wire  solvated_auto_mem_out_d_valid; // @[ComposerCore.scala 76:32]
  wire [3:0] solvated_auto_mem_out_d_bits_source; // @[ComposerCore.scala 76:32]
  wire  myWriters_WriteChannel_1_clock; // @[ComposerCore.scala 194:74]
  wire  myWriters_WriteChannel_1_reset; // @[ComposerCore.scala 194:74]
  wire  myWriters_WriteChannel_1_io_req_ready; // @[ComposerCore.scala 194:74]
  wire  myWriters_WriteChannel_1_io_req_valid; // @[ComposerCore.scala 194:74]
  wire [33:0] myWriters_WriteChannel_1_io_req_bits_addr; // @[ComposerCore.scala 194:74]
  wire [33:0] myWriters_WriteChannel_1_io_req_bits_len; // @[ComposerCore.scala 194:74]
  wire  myWriters_WriteChannel_1_io_channel_data_ready; // @[ComposerCore.scala 194:74]
  wire  myWriters_WriteChannel_1_io_channel_data_valid; // @[ComposerCore.scala 194:74]
  wire [31:0] myWriters_WriteChannel_1_io_channel_data_bits; // @[ComposerCore.scala 194:74]
  wire  myWriters_WriteChannel_1_io_channel_channelIdle; // @[ComposerCore.scala 194:74]
  wire  myWriters_WriteChannel_1_tl_out_a_ready; // @[ComposerCore.scala 194:74]
  wire  myWriters_WriteChannel_1_tl_out_a_valid; // @[ComposerCore.scala 194:74]
  wire  myWriters_WriteChannel_1_tl_out_a_bits_source; // @[ComposerCore.scala 194:74]
  wire [33:0] myWriters_WriteChannel_1_tl_out_a_bits_address; // @[ComposerCore.scala 194:74]
  wire [63:0] myWriters_WriteChannel_1_tl_out_a_bits_mask; // @[ComposerCore.scala 194:74]
  wire [511:0] myWriters_WriteChannel_1_tl_out_a_bits_data; // @[ComposerCore.scala 194:74]
  wire  myWriters_WriteChannel_1_tl_out_d_ready; // @[ComposerCore.scala 194:74]
  wire  myWriters_WriteChannel_1_tl_out_d_valid; // @[ComposerCore.scala 194:74]
  wire  myWriters_WriteChannel_1_tl_out_d_bits_source; // @[ComposerCore.scala 194:74]
  reg [2:0] state; // @[EnergyCalcTop.scala 31:22]
  reg [33:0] addr_data; // @[EnergyCalcTop.scala 32:52]
  reg [33:0] addr_HNBT; // @[EnergyCalcTop.scala 32:52]
  reg [31:0] sum; // @[EnergyCalcTop.scala 60:16]
  reg [31:0] a; // @[EnergyCalcTop.scala 61:23]
  reg [31:0] b; // @[EnergyCalcTop.scala 61:23]
  reg [31:0] c; // @[EnergyCalcTop.scala 61:23]
  reg [31:0] d; // @[EnergyCalcTop.scala 61:23]
  wire  _io_req_ready_T = state == 3'h0; // @[EnergyCalcTop.scala 64:25]
  wire  _T_1 = io_req_ready & io_req_valid; // @[Decoupled.scala 51:35]
  wire  _T_3 = ~reset; // @[EnergyCalcTop.scala 72:13]
  wire  _T_5 = io_req_bits_inst_rs1 == 5'h0; // @[EnergyCalcTop.scala 73:34]
  wire  _T_11 = io_req_bits_inst_rs1 == 5'h1; // @[EnergyCalcTop.scala 80:39]
  wire [2:0] _GEN_2 = io_req_bits_inst_rs1 == 5'h1 ? 3'h1 : state; // @[EnergyCalcTop.scala 80:83 84:15 31:22]
  wire  _T_14 = state == 3'h1; // @[EnergyCalcTop.scala 89:20]
  wire  _T_23 = state == 3'h2; // @[EnergyCalcTop.scala 113:20]
  wire [31:0] _GEN_18 = data_access_readReq_valid ? data_access_readRes_bits[31:0] : a; // @[EnergyCalcTop.scala 119:38 121:9 61:23]
  wire [31:0] _GEN_19 = data_access_readReq_valid ? data_access_readRes_bits[63:32] : b; // @[EnergyCalcTop.scala 119:38 122:9 61:23]
  wire [31:0] _GEN_20 = data_access_readReq_valid ? data_access_readRes_bits[95:64] : c; // @[EnergyCalcTop.scala 119:38 123:9 61:23]
  wire [31:0] _GEN_21 = data_access_readReq_valid ? data_access_readRes_bits[127:96] : d; // @[EnergyCalcTop.scala 119:38 124:9 61:23]
  wire [31:0] _sum_T_1 = a + b; // @[EnergyCalcTop.scala 130:14]
  wire [31:0] _sum_T_3 = _sum_T_1 + c; // @[EnergyCalcTop.scala 130:18]
  wire [31:0] _sum_T_5 = _sum_T_3 + d; // @[EnergyCalcTop.scala 130:22]
  wire  _T_30 = state == 3'h3; // @[EnergyCalcTop.scala 134:20]
  wire  _T_33 = myWriters_WriteChannel_1_io_channel_data_ready & myWriters_WriteChannel_1_io_channel_data_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_22 = _T_33 ? 3'h4 : state; // @[EnergyCalcTop.scala 138:30 140:13 31:22]
  wire  _T_36 = state == 3'h4; // @[EnergyCalcTop.scala 143:20]
  wire [2:0] _GEN_27 = myWriters_WriteChannel_1_io_channel_channelIdle ? 3'h5 : state; // @[EnergyCalcTop.scala 160:32 161:17 31:22]
  wire  _T_43 = state == 3'h5; // @[EnergyCalcTop.scala 164:20]
  wire  _T_46 = io_resp_ready & io_resp_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_28 = _T_46 ? 3'h0 : state; // @[EnergyCalcTop.scala 167:24 168:15 31:22]
  wire [2:0] _GEN_30 = state == 3'h5 ? _GEN_28 : state; // @[EnergyCalcTop.scala 164:34 31:22]
  wire [31:0] _GEN_33 = state == 3'h4 ? _GEN_18 : a; // @[EnergyCalcTop.scala 143:34 61:23]
  wire [31:0] _GEN_34 = state == 3'h4 ? _GEN_19 : b; // @[EnergyCalcTop.scala 143:34 61:23]
  wire [31:0] _GEN_35 = state == 3'h4 ? _GEN_20 : c; // @[EnergyCalcTop.scala 143:34 61:23]
  wire [31:0] _GEN_36 = state == 3'h4 ? _GEN_21 : d; // @[EnergyCalcTop.scala 143:34 61:23]
  wire [2:0] _GEN_37 = state == 3'h4 ? _GEN_27 : _GEN_30; // @[EnergyCalcTop.scala 143:34]
  wire  _GEN_38 = state == 3'h4 ? 1'h0 : _T_43; // @[EnergyCalcTop.scala 143:34 65:17]
  wire [2:0] _GEN_40 = state == 3'h3 ? _GEN_22 : _GEN_37; // @[EnergyCalcTop.scala 134:33]
  wire  _GEN_47 = state == 3'h3 ? 1'h0 : _GEN_38; // @[EnergyCalcTop.scala 134:33 65:17]
  wire  _GEN_48 = state == 3'h2 ? state == 3'h2 : _T_36; // @[EnergyCalcTop.scala 113:37 115:31]
  wire  _GEN_56 = state == 3'h2 ? 1'h0 : _T_30; // @[EnergyCalcTop.scala 113:37 62:23]
  wire  _GEN_57 = state == 3'h2 ? 1'h0 : _GEN_47; // @[EnergyCalcTop.scala 113:37 65:17]
  wire  _GEN_66 = state == 3'h1 ? 1'h0 : _GEN_56; // @[EnergyCalcTop.scala 62:23 89:32]
  wire  _GEN_67 = state == 3'h1 ? 1'h0 : _GEN_57; // @[EnergyCalcTop.scala 65:17 89:32]
  wire  _GEN_82 = _io_req_ready_T & _T_1; // @[EnergyCalcTop.scala 72:13]
  wire  _GEN_84 = _GEN_82 & _T_5; // @[EnergyCalcTop.scala 77:15]
  wire  _GEN_91 = ~_io_req_ready_T; // @[EnergyCalcTop.scala 90:11]
  wire  _GEN_92 = ~_io_req_ready_T & _T_14; // @[EnergyCalcTop.scala 90:11]
  wire  _GEN_97 = _GEN_92 & data_access_readRes_valid; // @[EnergyCalcTop.scala 101:13]
  wire  _GEN_103 = _GEN_91 & ~_T_14; // @[EnergyCalcTop.scala 114:11]
  wire  _GEN_104 = _GEN_91 & ~_T_14 & _T_23; // @[EnergyCalcTop.scala 114:11]
  wire  _GEN_118 = _GEN_103 & ~_T_23; // @[EnergyCalcTop.scala 135:11]
  wire  _GEN_119 = _GEN_103 & ~_T_23 & _T_30; // @[EnergyCalcTop.scala 135:11]
  wire  _GEN_133 = _GEN_118 & ~_T_30; // @[EnergyCalcTop.scala 154:13]
  wire  _GEN_134 = _GEN_118 & ~_T_30 & _T_36; // @[EnergyCalcTop.scala 154:13]
  CScratchpad data ( // @[ComposerCore.scala 76:32]
    .clock(data_clock),
    .reset(data_reset),
    .auto_mem_out_a_ready(data_auto_mem_out_a_ready),
    .auto_mem_out_a_valid(data_auto_mem_out_a_valid),
    .auto_mem_out_a_bits_size(data_auto_mem_out_a_bits_size),
    .auto_mem_out_a_bits_source(data_auto_mem_out_a_bits_source),
    .auto_mem_out_a_bits_address(data_auto_mem_out_a_bits_address),
    .auto_mem_out_a_bits_mask(data_auto_mem_out_a_bits_mask),
    .auto_mem_out_d_ready(data_auto_mem_out_d_ready),
    .auto_mem_out_d_valid(data_auto_mem_out_d_valid),
    .auto_mem_out_d_bits_source(data_auto_mem_out_d_bits_source),
    .auto_mem_out_d_bits_data(data_auto_mem_out_d_bits_data),
    .access_readReq_valid(data_access_readReq_valid),
    .access_readRes_valid(data_access_readRes_valid),
    .access_readRes_bits(data_access_readRes_bits)
  );
  CScratchpad_1 halfNonBonded ( // @[ComposerCore.scala 76:32]
    .clock(halfNonBonded_clock),
    .reset(halfNonBonded_reset),
    .auto_mem_out_a_ready(halfNonBonded_auto_mem_out_a_ready),
    .auto_mem_out_a_valid(halfNonBonded_auto_mem_out_a_valid),
    .auto_mem_out_a_bits_size(halfNonBonded_auto_mem_out_a_bits_size),
    .auto_mem_out_a_bits_source(halfNonBonded_auto_mem_out_a_bits_source),
    .auto_mem_out_a_bits_address(halfNonBonded_auto_mem_out_a_bits_address),
    .auto_mem_out_a_bits_mask(halfNonBonded_auto_mem_out_a_bits_mask),
    .auto_mem_out_d_ready(halfNonBonded_auto_mem_out_d_ready),
    .auto_mem_out_d_valid(halfNonBonded_auto_mem_out_d_valid),
    .auto_mem_out_d_bits_source(halfNonBonded_auto_mem_out_d_bits_source)
  );
  CScratchpad_2 nonBonded ( // @[ComposerCore.scala 76:32]
    .clock(nonBonded_clock),
    .reset(nonBonded_reset),
    .auto_mem_out_a_ready(nonBonded_auto_mem_out_a_ready),
    .auto_mem_out_a_valid(nonBonded_auto_mem_out_a_valid),
    .auto_mem_out_a_bits_size(nonBonded_auto_mem_out_a_bits_size),
    .auto_mem_out_a_bits_source(nonBonded_auto_mem_out_a_bits_source),
    .auto_mem_out_a_bits_address(nonBonded_auto_mem_out_a_bits_address),
    .auto_mem_out_a_bits_mask(nonBonded_auto_mem_out_a_bits_mask),
    .auto_mem_out_d_ready(nonBonded_auto_mem_out_d_ready),
    .auto_mem_out_d_valid(nonBonded_auto_mem_out_d_valid),
    .auto_mem_out_d_bits_source(nonBonded_auto_mem_out_d_bits_source)
  );
  CScratchpad_3 solvated ( // @[ComposerCore.scala 76:32]
    .clock(solvated_clock),
    .reset(solvated_reset),
    .auto_mem_out_a_ready(solvated_auto_mem_out_a_ready),
    .auto_mem_out_a_valid(solvated_auto_mem_out_a_valid),
    .auto_mem_out_a_bits_size(solvated_auto_mem_out_a_bits_size),
    .auto_mem_out_a_bits_source(solvated_auto_mem_out_a_bits_source),
    .auto_mem_out_a_bits_address(solvated_auto_mem_out_a_bits_address),
    .auto_mem_out_a_bits_mask(solvated_auto_mem_out_a_bits_mask),
    .auto_mem_out_d_ready(solvated_auto_mem_out_d_ready),
    .auto_mem_out_d_valid(solvated_auto_mem_out_d_valid),
    .auto_mem_out_d_bits_source(solvated_auto_mem_out_d_bits_source)
  );
  SequentialWriter myWriters_WriteChannel_1 ( // @[ComposerCore.scala 194:74]
    .clock(myWriters_WriteChannel_1_clock),
    .reset(myWriters_WriteChannel_1_reset),
    .io_req_ready(myWriters_WriteChannel_1_io_req_ready),
    .io_req_valid(myWriters_WriteChannel_1_io_req_valid),
    .io_req_bits_addr(myWriters_WriteChannel_1_io_req_bits_addr),
    .io_req_bits_len(myWriters_WriteChannel_1_io_req_bits_len),
    .io_channel_data_ready(myWriters_WriteChannel_1_io_channel_data_ready),
    .io_channel_data_valid(myWriters_WriteChannel_1_io_channel_data_valid),
    .io_channel_data_bits(myWriters_WriteChannel_1_io_channel_data_bits),
    .io_channel_channelIdle(myWriters_WriteChannel_1_io_channel_channelIdle),
    .tl_out_a_ready(myWriters_WriteChannel_1_tl_out_a_ready),
    .tl_out_a_valid(myWriters_WriteChannel_1_tl_out_a_valid),
    .tl_out_a_bits_source(myWriters_WriteChannel_1_tl_out_a_bits_source),
    .tl_out_a_bits_address(myWriters_WriteChannel_1_tl_out_a_bits_address),
    .tl_out_a_bits_mask(myWriters_WriteChannel_1_tl_out_a_bits_mask),
    .tl_out_a_bits_data(myWriters_WriteChannel_1_tl_out_a_bits_data),
    .tl_out_d_ready(myWriters_WriteChannel_1_tl_out_d_ready),
    .tl_out_d_valid(myWriters_WriteChannel_1_tl_out_d_valid),
    .tl_out_d_bits_source(myWriters_WriteChannel_1_tl_out_d_bits_source)
  );
  assign auto_solvated_mem_out_a_valid = solvated_auto_mem_out_a_valid; // @[LazyModule.scala 368:12]
  assign auto_solvated_mem_out_a_bits_size = solvated_auto_mem_out_a_bits_size; // @[LazyModule.scala 368:12]
  assign auto_solvated_mem_out_a_bits_source = solvated_auto_mem_out_a_bits_source; // @[LazyModule.scala 368:12]
  assign auto_solvated_mem_out_a_bits_address = solvated_auto_mem_out_a_bits_address; // @[LazyModule.scala 368:12]
  assign auto_solvated_mem_out_a_bits_mask = solvated_auto_mem_out_a_bits_mask; // @[LazyModule.scala 368:12]
  assign auto_solvated_mem_out_d_ready = solvated_auto_mem_out_d_ready; // @[LazyModule.scala 368:12]
  assign auto_nonBonded_mem_out_a_valid = nonBonded_auto_mem_out_a_valid; // @[LazyModule.scala 368:12]
  assign auto_nonBonded_mem_out_a_bits_size = nonBonded_auto_mem_out_a_bits_size; // @[LazyModule.scala 368:12]
  assign auto_nonBonded_mem_out_a_bits_source = nonBonded_auto_mem_out_a_bits_source; // @[LazyModule.scala 368:12]
  assign auto_nonBonded_mem_out_a_bits_address = nonBonded_auto_mem_out_a_bits_address; // @[LazyModule.scala 368:12]
  assign auto_nonBonded_mem_out_a_bits_mask = nonBonded_auto_mem_out_a_bits_mask; // @[LazyModule.scala 368:12]
  assign auto_nonBonded_mem_out_d_ready = nonBonded_auto_mem_out_d_ready; // @[LazyModule.scala 368:12]
  assign auto_halfNonBonded_mem_out_a_valid = halfNonBonded_auto_mem_out_a_valid; // @[LazyModule.scala 368:12]
  assign auto_halfNonBonded_mem_out_a_bits_size = halfNonBonded_auto_mem_out_a_bits_size; // @[LazyModule.scala 368:12]
  assign auto_halfNonBonded_mem_out_a_bits_source = halfNonBonded_auto_mem_out_a_bits_source; // @[LazyModule.scala 368:12]
  assign auto_halfNonBonded_mem_out_a_bits_address = halfNonBonded_auto_mem_out_a_bits_address; // @[LazyModule.scala 368:12]
  assign auto_halfNonBonded_mem_out_a_bits_mask = halfNonBonded_auto_mem_out_a_bits_mask; // @[LazyModule.scala 368:12]
  assign auto_halfNonBonded_mem_out_d_ready = halfNonBonded_auto_mem_out_d_ready; // @[LazyModule.scala 368:12]
  assign auto_data_mem_out_a_valid = data_auto_mem_out_a_valid; // @[LazyModule.scala 368:12]
  assign auto_data_mem_out_a_bits_size = data_auto_mem_out_a_bits_size; // @[LazyModule.scala 368:12]
  assign auto_data_mem_out_a_bits_source = data_auto_mem_out_a_bits_source; // @[LazyModule.scala 368:12]
  assign auto_data_mem_out_a_bits_address = data_auto_mem_out_a_bits_address; // @[LazyModule.scala 368:12]
  assign auto_data_mem_out_a_bits_mask = data_auto_mem_out_a_bits_mask; // @[LazyModule.scala 368:12]
  assign auto_data_mem_out_d_ready = data_auto_mem_out_d_ready; // @[LazyModule.scala 368:12]
  assign auto_writers_out_a_valid = myWriters_WriteChannel_1_tl_out_a_valid; // @[Nodes.scala 1212:84 ComposerCore.scala 198:16]
  assign auto_writers_out_a_bits_source = myWriters_WriteChannel_1_tl_out_a_bits_source; // @[Nodes.scala 1212:84 ComposerCore.scala 198:16]
  assign auto_writers_out_a_bits_address = myWriters_WriteChannel_1_tl_out_a_bits_address; // @[Nodes.scala 1212:84 ComposerCore.scala 198:16]
  assign auto_writers_out_a_bits_mask = myWriters_WriteChannel_1_tl_out_a_bits_mask; // @[Nodes.scala 1212:84 ComposerCore.scala 198:16]
  assign auto_writers_out_a_bits_data = myWriters_WriteChannel_1_tl_out_a_bits_data; // @[Nodes.scala 1212:84 ComposerCore.scala 198:16]
  assign auto_writers_out_d_ready = myWriters_WriteChannel_1_tl_out_d_ready; // @[Nodes.scala 1212:84 ComposerCore.scala 198:16]
  assign io_req_ready = state == 3'h0; // @[EnergyCalcTop.scala 64:25]
  assign io_resp_valid = _io_req_ready_T ? 1'h0 : _GEN_67; // @[EnergyCalcTop.scala 65:17 70:27]
  assign data_clock = clock;
  assign data_reset = reset;
  assign data_auto_mem_out_a_ready = auto_data_mem_out_a_ready; // @[LazyModule.scala 368:12]
  assign data_auto_mem_out_d_valid = auto_data_mem_out_d_valid; // @[LazyModule.scala 368:12]
  assign data_auto_mem_out_d_bits_source = auto_data_mem_out_d_bits_source; // @[LazyModule.scala 368:12]
  assign data_auto_mem_out_d_bits_data = auto_data_mem_out_d_bits_data; // @[LazyModule.scala 368:12]
  assign data_access_readReq_valid = state == 3'h1 ? state == 3'h1 : _GEN_48; // @[EnergyCalcTop.scala 89:32 91:31]
  assign halfNonBonded_clock = clock;
  assign halfNonBonded_reset = reset;
  assign halfNonBonded_auto_mem_out_a_ready = auto_halfNonBonded_mem_out_a_ready; // @[LazyModule.scala 368:12]
  assign halfNonBonded_auto_mem_out_d_valid = auto_halfNonBonded_mem_out_d_valid; // @[LazyModule.scala 368:12]
  assign halfNonBonded_auto_mem_out_d_bits_source = auto_halfNonBonded_mem_out_d_bits_source; // @[LazyModule.scala 368:12]
  assign nonBonded_clock = clock;
  assign nonBonded_reset = reset;
  assign nonBonded_auto_mem_out_a_ready = auto_nonBonded_mem_out_a_ready; // @[LazyModule.scala 368:12]
  assign nonBonded_auto_mem_out_d_valid = auto_nonBonded_mem_out_d_valid; // @[LazyModule.scala 368:12]
  assign nonBonded_auto_mem_out_d_bits_source = auto_nonBonded_mem_out_d_bits_source; // @[LazyModule.scala 368:12]
  assign solvated_clock = clock;
  assign solvated_reset = reset;
  assign solvated_auto_mem_out_a_ready = auto_solvated_mem_out_a_ready; // @[LazyModule.scala 368:12]
  assign solvated_auto_mem_out_d_valid = auto_solvated_mem_out_d_valid; // @[LazyModule.scala 368:12]
  assign solvated_auto_mem_out_d_bits_source = auto_solvated_mem_out_d_bits_source; // @[LazyModule.scala 368:12]
  assign myWriters_WriteChannel_1_clock = clock;
  assign myWriters_WriteChannel_1_reset = reset;
  assign myWriters_WriteChannel_1_io_req_valid = myWriters_WriteChannel_valid; // @[ComposerCore.scala 202:15]
  assign myWriters_WriteChannel_1_io_req_bits_addr = myWriters_WriteChannel_bits_addr; // @[ComposerCore.scala 202:15]
  assign myWriters_WriteChannel_1_io_req_bits_len = myWriters_WriteChannel_bits_len; // @[ComposerCore.scala 202:15]
  assign myWriters_WriteChannel_1_io_channel_data_valid = _io_req_ready_T ? 1'h0 : _GEN_66; // @[EnergyCalcTop.scala 62:23 70:27]
  assign myWriters_WriteChannel_1_io_channel_data_bits = sum; // @[EnergyCalcTop.scala 63:22]
  assign myWriters_WriteChannel_1_tl_out_a_ready = auto_writers_out_a_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign myWriters_WriteChannel_1_tl_out_d_valid = auto_writers_out_d_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign myWriters_WriteChannel_1_tl_out_d_bits_source = auto_writers_out_d_bits_source; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  always @(posedge clock) begin
    if (reset) begin // @[EnergyCalcTop.scala 31:22]
      state <= 3'h0; // @[EnergyCalcTop.scala 31:22]
    end else if (_io_req_ready_T) begin // @[EnergyCalcTop.scala 70:27]
      if (_T_1) begin // @[EnergyCalcTop.scala 71:23]
        if (!(io_req_bits_inst_rs1 == 5'h0)) begin // @[EnergyCalcTop.scala 73:81]
          state <= _GEN_2;
        end
      end
    end else if (state == 3'h1) begin // @[EnergyCalcTop.scala 89:32]
      if (data_access_readRes_valid) begin // @[EnergyCalcTop.scala 95:38]
        state <= 3'h2; // @[EnergyCalcTop.scala 105:13]
      end
    end else if (state == 3'h2) begin // @[EnergyCalcTop.scala 113:37]
      state <= 3'h3; // @[EnergyCalcTop.scala 132:11]
    end else begin
      state <= _GEN_40;
    end
    if (_io_req_ready_T) begin // @[EnergyCalcTop.scala 70:27]
      if (_T_1) begin // @[EnergyCalcTop.scala 71:23]
        if (io_req_bits_inst_rs1 == 5'h0) begin // @[EnergyCalcTop.scala 73:81]
          addr_data <= io_req_bits_payload1[33:0]; // @[EnergyCalcTop.scala 74:19]
        end
      end
    end
    if (_io_req_ready_T) begin // @[EnergyCalcTop.scala 70:27]
      if (_T_1) begin // @[EnergyCalcTop.scala 71:23]
        if (io_req_bits_inst_rs1 == 5'h0) begin // @[EnergyCalcTop.scala 73:81]
          addr_HNBT <= io_req_bits_payload2[33:0]; // @[EnergyCalcTop.scala 75:19]
        end
      end
    end
    if (!(_io_req_ready_T)) begin // @[EnergyCalcTop.scala 70:27]
      if (!(state == 3'h1)) begin // @[EnergyCalcTop.scala 89:32]
        if (state == 3'h2) begin // @[EnergyCalcTop.scala 113:37]
          sum <= _sum_T_5; // @[EnergyCalcTop.scala 130:9]
        end
      end
    end
    if (!(_io_req_ready_T)) begin // @[EnergyCalcTop.scala 70:27]
      if (state == 3'h1) begin // @[EnergyCalcTop.scala 89:32]
        if (data_access_readRes_valid) begin // @[EnergyCalcTop.scala 95:38]
          a <= data_access_readRes_bits[31:0]; // @[EnergyCalcTop.scala 97:9]
        end
      end else if (state == 3'h2) begin // @[EnergyCalcTop.scala 113:37]
        if (data_access_readReq_valid) begin // @[EnergyCalcTop.scala 119:38]
          a <= data_access_readRes_bits[31:0]; // @[EnergyCalcTop.scala 121:9]
        end
      end else if (!(state == 3'h3)) begin // @[EnergyCalcTop.scala 134:33]
        a <= _GEN_33;
      end
    end
    if (!(_io_req_ready_T)) begin // @[EnergyCalcTop.scala 70:27]
      if (state == 3'h1) begin // @[EnergyCalcTop.scala 89:32]
        if (data_access_readRes_valid) begin // @[EnergyCalcTop.scala 95:38]
          b <= data_access_readRes_bits[63:32]; // @[EnergyCalcTop.scala 98:9]
        end
      end else if (state == 3'h2) begin // @[EnergyCalcTop.scala 113:37]
        if (data_access_readReq_valid) begin // @[EnergyCalcTop.scala 119:38]
          b <= data_access_readRes_bits[63:32]; // @[EnergyCalcTop.scala 122:9]
        end
      end else if (!(state == 3'h3)) begin // @[EnergyCalcTop.scala 134:33]
        b <= _GEN_34;
      end
    end
    if (!(_io_req_ready_T)) begin // @[EnergyCalcTop.scala 70:27]
      if (state == 3'h1) begin // @[EnergyCalcTop.scala 89:32]
        if (data_access_readRes_valid) begin // @[EnergyCalcTop.scala 95:38]
          c <= data_access_readRes_bits[95:64]; // @[EnergyCalcTop.scala 99:9]
        end
      end else if (state == 3'h2) begin // @[EnergyCalcTop.scala 113:37]
        if (data_access_readReq_valid) begin // @[EnergyCalcTop.scala 119:38]
          c <= data_access_readRes_bits[95:64]; // @[EnergyCalcTop.scala 123:9]
        end
      end else if (!(state == 3'h3)) begin // @[EnergyCalcTop.scala 134:33]
        c <= _GEN_35;
      end
    end
    if (!(_io_req_ready_T)) begin // @[EnergyCalcTop.scala 70:27]
      if (state == 3'h1) begin // @[EnergyCalcTop.scala 89:32]
        if (data_access_readRes_valid) begin // @[EnergyCalcTop.scala 95:38]
          d <= data_access_readRes_bits[127:96]; // @[EnergyCalcTop.scala 100:9]
        end
      end else if (state == 3'h2) begin // @[EnergyCalcTop.scala 113:37]
        if (data_access_readReq_valid) begin // @[EnergyCalcTop.scala 119:38]
          d <= data_access_readRes_bits[127:96]; // @[EnergyCalcTop.scala 124:9]
        end
      end else if (!(state == 3'h3)) begin // @[EnergyCalcTop.scala 134:33]
        d <= _GEN_36;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_io_req_ready_T & _T_1 & ~reset) begin
          $fwrite(32'h80000002,"input fired\n"); // @[EnergyCalcTop.scala 72:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_82 & _T_5 & _T_3) begin
          $fwrite(32'h80000002,"input 1 data address %b\n",addr_data); // @[EnergyCalcTop.scala 77:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_84 & _T_3) begin
          $fwrite(32'h80000002,"input 1 HNBT address %d\n",addr_HNBT); // @[EnergyCalcTop.scala 78:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_82 & ~_T_5 & _T_11 & _T_3) begin
          $fwrite(32'h80000002,"input 2\n"); // @[EnergyCalcTop.scala 83:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_io_req_ready_T & _T_14 & _T_3) begin
          $fwrite(32'h80000002,"read\n"); // @[EnergyCalcTop.scala 90:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_92 & _T_3) begin
          $fwrite(32'h80000002,"input 1 data address %b\n",addr_HNBT); // @[EnergyCalcTop.scala 94:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_92 & data_access_readRes_valid & _T_3) begin
          $fwrite(32'h80000002,"%b\n",data_access_readRes_bits); // @[EnergyCalcTop.scala 101:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_97 & _T_3) begin
          $fwrite(32'h80000002,"a%d b%d c%d d%d\n",a,b,c,d); // @[EnergyCalcTop.scala 103:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_91 & ~_T_14 & _T_23 & _T_3) begin
          $fwrite(32'h80000002,"calculate\n"); // @[EnergyCalcTop.scala 114:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_104 & data_access_readReq_valid & _T_3) begin
          $fwrite(32'h80000002,"%b\n",data_access_readRes_bits); // @[EnergyCalcTop.scala 125:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_104 & _T_3) begin
          $fwrite(32'h80000002,"a%d b%d c%d d%d\n",a,b,c,d); // @[EnergyCalcTop.scala 128:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & ~_T_23 & _T_30 & _T_3) begin
          $fwrite(32'h80000002,"store\n"); // @[EnergyCalcTop.scala 135:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_119 & _T_33 & _T_3) begin
          $fwrite(32'h80000002,"output sum - %d\n",sum); // @[EnergyCalcTop.scala 139:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_118 & ~_T_30 & _T_36 & data_access_readReq_valid & _T_3) begin
          $fwrite(32'h80000002,"%b\n",data_access_readRes_bits); // @[EnergyCalcTop.scala 154:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_134 & _T_3) begin
          $fwrite(32'h80000002,"a%d b%d c%d d%d\n",a,b,c,d); // @[EnergyCalcTop.scala 157:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_134 & _T_3) begin
          $fwrite(32'h80000002,"commit\n"); // @[EnergyCalcTop.scala 159:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & ~_T_36 & _T_43 & _T_3) begin
          $fwrite(32'h80000002,"finish\n"); // @[EnergyCalcTop.scala 165:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module MultiLevelArbiter(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [59:0] io_in_0_bits_data,
  input  [4:0]  io_in_0_bits_rd,
  input         io_out_ready,
  output        io_out_valid,
  output [59:0] io_out_bits_data,
  output [4:0]  io_out_bits_rd
);
  assign io_in_0_ready = io_out_ready; // @[MultiLevelArbiter.scala 55:14]
  assign io_out_valid = io_in_0_valid; // @[MultiLevelArbiter.scala 55:14]
  assign io_out_bits_data = io_in_0_bits_data; // @[MultiLevelArbiter.scala 55:14]
  assign io_out_bits_rd = io_in_0_bits_rd; // @[MultiLevelArbiter.scala 55:14]
endmodule
module RRArbiter(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [4:0]  io_in_0_bits_inst_rs1,
  input  [4:0]  io_in_0_bits_inst_rs2,
  input  [2:0]  io_in_0_bits_inst_funct,
  input  [7:0]  io_in_0_bits_core_id,
  input  [55:0] io_in_0_bits_payload1,
  input  [63:0] io_in_0_bits_payload2,
  input         io_out_ready,
  output        io_out_valid,
  output [4:0]  io_out_bits_inst_rs1,
  output [4:0]  io_out_bits_inst_rs2,
  output [2:0]  io_out_bits_inst_funct,
  output [7:0]  io_out_bits_core_id,
  output [55:0] io_out_bits_payload1,
  output [63:0] io_out_bits_payload2
);
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 74:21]
  assign io_out_valid = io_in_0_valid; // @[Arbiter.scala 55:16]
  assign io_out_bits_inst_rs1 = io_in_0_bits_inst_rs1; // @[Arbiter.scala 56:15]
  assign io_out_bits_inst_rs2 = io_in_0_bits_inst_rs2; // @[Arbiter.scala 56:15]
  assign io_out_bits_inst_funct = io_in_0_bits_inst_funct; // @[Arbiter.scala 56:15]
  assign io_out_bits_core_id = io_in_0_bits_core_id; // @[Arbiter.scala 56:15]
  assign io_out_bits_payload1 = io_in_0_bits_payload1; // @[Arbiter.scala 56:15]
  assign io_out_bits_payload2 = io_in_0_bits_payload2; // @[Arbiter.scala 56:15]
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [4:0]  io_enq_bits_inst_rs1,
  input  [4:0]  io_enq_bits_inst_rs2,
  input  [2:0]  io_enq_bits_inst_funct,
  input  [7:0]  io_enq_bits_core_id,
  input  [55:0] io_enq_bits_payload1,
  input  [63:0] io_enq_bits_payload2,
  input         io_deq_ready,
  output        io_deq_valid,
  output [4:0]  io_deq_bits_inst_rs1,
  output [4:0]  io_deq_bits_inst_rs2,
  output [2:0]  io_deq_bits_inst_funct,
  output [7:0]  io_deq_bits_core_id,
  output [55:0] io_deq_bits_payload1,
  output [63:0] io_deq_bits_payload2
);
  reg [4:0] ram_inst_rs1 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_inst_rs1_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_inst_rs1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [4:0] ram_inst_rs1_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [4:0] ram_inst_rs1_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_inst_rs1_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_inst_rs1_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_inst_rs1_MPORT_en; // @[Decoupled.scala 273:95]
  reg [4:0] ram_inst_rs2 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_inst_rs2_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_inst_rs2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [4:0] ram_inst_rs2_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [4:0] ram_inst_rs2_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_inst_rs2_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_inst_rs2_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_inst_rs2_MPORT_en; // @[Decoupled.scala 273:95]
  reg [2:0] ram_inst_funct [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_inst_funct_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_inst_funct_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [2:0] ram_inst_funct_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_inst_funct_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_inst_funct_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_inst_funct_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_inst_funct_MPORT_en; // @[Decoupled.scala 273:95]
  reg [7:0] ram_core_id [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_core_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_core_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [7:0] ram_core_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [7:0] ram_core_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_core_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_core_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_core_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [55:0] ram_payload1 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_payload1_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_payload1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [55:0] ram_payload1_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [55:0] ram_payload1_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_payload1_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_payload1_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_payload1_MPORT_en; // @[Decoupled.scala 273:95]
  reg [63:0] ram_payload2 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_payload2_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_payload2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload2_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload2_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_payload2_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_payload2_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_payload2_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_inst_rs1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_inst_rs1_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_inst_rs1_io_deq_bits_MPORT_data = ram_inst_rs1[ram_inst_rs1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_inst_rs1_MPORT_data = io_enq_bits_inst_rs1;
  assign ram_inst_rs1_MPORT_addr = enq_ptr_value;
  assign ram_inst_rs1_MPORT_mask = 1'h1;
  assign ram_inst_rs1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_inst_rs2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_inst_rs2_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_inst_rs2_io_deq_bits_MPORT_data = ram_inst_rs2[ram_inst_rs2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_inst_rs2_MPORT_data = io_enq_bits_inst_rs2;
  assign ram_inst_rs2_MPORT_addr = enq_ptr_value;
  assign ram_inst_rs2_MPORT_mask = 1'h1;
  assign ram_inst_rs2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_inst_funct_io_deq_bits_MPORT_en = 1'h1;
  assign ram_inst_funct_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_inst_funct_io_deq_bits_MPORT_data = ram_inst_funct[ram_inst_funct_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_inst_funct_MPORT_data = io_enq_bits_inst_funct;
  assign ram_inst_funct_MPORT_addr = enq_ptr_value;
  assign ram_inst_funct_MPORT_mask = 1'h1;
  assign ram_inst_funct_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_core_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_core_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_core_id_io_deq_bits_MPORT_data = ram_core_id[ram_core_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_core_id_MPORT_data = io_enq_bits_core_id;
  assign ram_core_id_MPORT_addr = enq_ptr_value;
  assign ram_core_id_MPORT_mask = 1'h1;
  assign ram_core_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_payload1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_payload1_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_payload1_io_deq_bits_MPORT_data = ram_payload1[ram_payload1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_payload1_MPORT_data = io_enq_bits_payload1;
  assign ram_payload1_MPORT_addr = enq_ptr_value;
  assign ram_payload1_MPORT_mask = 1'h1;
  assign ram_payload1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_payload2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_payload2_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_payload2_io_deq_bits_MPORT_data = ram_payload2[ram_payload2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_payload2_MPORT_data = io_enq_bits_payload2;
  assign ram_payload2_MPORT_addr = enq_ptr_value;
  assign ram_payload2_MPORT_mask = 1'h1;
  assign ram_payload2_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_inst_rs1 = ram_inst_rs1_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_inst_rs2 = ram_inst_rs2_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_inst_funct = ram_inst_funct_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_core_id = ram_core_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_payload1 = ram_payload1_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_payload2 = ram_payload2_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_inst_rs1_MPORT_en & ram_inst_rs1_MPORT_mask) begin
      ram_inst_rs1[ram_inst_rs1_MPORT_addr] <= ram_inst_rs1_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_inst_rs2_MPORT_en & ram_inst_rs2_MPORT_mask) begin
      ram_inst_rs2[ram_inst_rs2_MPORT_addr] <= ram_inst_rs2_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_inst_funct_MPORT_en & ram_inst_funct_MPORT_mask) begin
      ram_inst_funct[ram_inst_funct_MPORT_addr] <= ram_inst_funct_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_core_id_MPORT_en & ram_core_id_MPORT_mask) begin
      ram_core_id[ram_core_id_MPORT_addr] <= ram_core_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_payload1_MPORT_en & ram_payload1_MPORT_mask) begin
      ram_payload1[ram_payload1_MPORT_addr] <= ram_payload1_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_payload2_MPORT_en & ram_payload2_MPORT_mask) begin
      ram_payload2[ram_payload2_MPORT_addr] <= ram_payload2_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
endmodule
module Queue_1(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_deq_ready,
  output        io_deq_valid,
  output [59:0] io_deq_bits_data,
  output [4:0]  io_deq_bits_rd
);
  reg [59:0] ram_data [0:3]; // @[Decoupled.scala 273:44]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [1:0] ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire [59:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire [59:0] ram_data_MPORT_data; // @[Decoupled.scala 273:44]
  wire [1:0] ram_data_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_data_io_deq_bits_MPORT_en_pipe_0;
  reg [1:0] ram_data_io_deq_bits_MPORT_addr_pipe_0;
  reg [4:0] ram_rd [0:3]; // @[Decoupled.scala 273:44]
  wire  ram_rd_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [1:0] ram_rd_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire [4:0] ram_rd_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire [4:0] ram_rd_MPORT_data; // @[Decoupled.scala 273:44]
  wire [1:0] ram_rd_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_rd_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_rd_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_rd_io_deq_bits_MPORT_en_pipe_0;
  reg [1:0] ram_rd_io_deq_bits_MPORT_addr_pipe_0;
  reg [1:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire [2:0] _deq_ptr_next_T_1 = 3'h4 - 3'h1; // @[Decoupled.scala 306:57]
  wire [2:0] _GEN_16 = {{1'd0}, deq_ptr_value}; // @[Decoupled.scala 306:42]
  assign ram_data_io_deq_bits_MPORT_en = ram_data_io_deq_bits_MPORT_en_pipe_0;
  assign ram_data_io_deq_bits_MPORT_addr = ram_data_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_data_MPORT_data = 60'h0;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_rd_io_deq_bits_MPORT_en = ram_rd_io_deq_bits_MPORT_en_pipe_0;
  assign ram_rd_io_deq_bits_MPORT_addr = ram_rd_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_rd_io_deq_bits_MPORT_data = ram_rd[ram_rd_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_rd_MPORT_data = 5'h0;
  assign ram_rd_MPORT_addr = enq_ptr_value;
  assign ram_rd_MPORT_mask = 1'h1;
  assign ram_rd_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_rd = ram_rd_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  always @(posedge clock) begin
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_data_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_16 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_data_io_deq_bits_MPORT_addr_pipe_0 <= 2'h0;
        end else begin
          ram_data_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_data_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_rd_MPORT_en & ram_rd_MPORT_mask) begin
      ram_rd[ram_rd_MPORT_addr] <= ram_rd_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_rd_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_16 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_rd_io_deq_bits_MPORT_addr_pipe_0 <= 2'h0;
        end else begin
          ram_rd_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_rd_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
endmodule
module Queue_2(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [4:0]  io_enq_bits_rd,
  input  [46:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [4:0]  io_deq_bits_rd,
  output [3:0]  io_deq_bits_system_id,
  output [7:0]  io_deq_bits_core_id,
  output [46:0] io_deq_bits_data
);
  reg [4:0] ram_rd [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_rd_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_rd_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [4:0] ram_rd_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [4:0] ram_rd_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_rd_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_rd_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_rd_MPORT_en; // @[Decoupled.scala 273:95]
  reg [3:0] ram_system_id [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_system_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_system_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [3:0] ram_system_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [3:0] ram_system_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_system_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_system_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_system_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [7:0] ram_core_id [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_core_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_core_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [7:0] ram_core_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [7:0] ram_core_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_core_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_core_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_core_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [46:0] ram_data [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [46:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [46:0] ram_data_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_rd_io_deq_bits_MPORT_en = 1'h1;
  assign ram_rd_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_rd_io_deq_bits_MPORT_data = ram_rd[ram_rd_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_rd_MPORT_data = io_enq_bits_rd;
  assign ram_rd_MPORT_addr = enq_ptr_value;
  assign ram_rd_MPORT_mask = 1'h1;
  assign ram_rd_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_system_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_system_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_system_id_io_deq_bits_MPORT_data = ram_system_id[ram_system_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_system_id_MPORT_data = 4'h0;
  assign ram_system_id_MPORT_addr = enq_ptr_value;
  assign ram_system_id_MPORT_mask = 1'h1;
  assign ram_system_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_core_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_core_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_core_id_io_deq_bits_MPORT_data = ram_core_id[ram_core_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_core_id_MPORT_data = 8'h0;
  assign ram_core_id_MPORT_addr = enq_ptr_value;
  assign ram_core_id_MPORT_mask = 1'h1;
  assign ram_core_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_rd = ram_rd_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_system_id = ram_system_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_core_id = ram_core_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_rd_MPORT_en & ram_rd_MPORT_mask) begin
      ram_rd[ram_rd_MPORT_addr] <= ram_rd_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_system_id_MPORT_en & ram_system_id_MPORT_mask) begin
      ram_system_id[ram_system_id_MPORT_addr] <= ram_system_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_core_id_MPORT_en & ram_core_id_MPORT_mask) begin
      ram_core_id[ram_core_id_MPORT_addr] <= ram_core_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
endmodule
module ComposerSystem(
  input          clock,
  input          reset,
  input          auto_memory_endpoint_identity_out_4_a_ready,
  output         auto_memory_endpoint_identity_out_4_a_valid,
  output [2:0]   auto_memory_endpoint_identity_out_4_a_bits_size,
  output [3:0]   auto_memory_endpoint_identity_out_4_a_bits_source,
  output [33:0]  auto_memory_endpoint_identity_out_4_a_bits_address,
  output [63:0]  auto_memory_endpoint_identity_out_4_a_bits_mask,
  output         auto_memory_endpoint_identity_out_4_d_ready,
  input          auto_memory_endpoint_identity_out_4_d_valid,
  input  [3:0]   auto_memory_endpoint_identity_out_4_d_bits_source,
  input          auto_memory_endpoint_identity_out_3_a_ready,
  output         auto_memory_endpoint_identity_out_3_a_valid,
  output [2:0]   auto_memory_endpoint_identity_out_3_a_bits_size,
  output [3:0]   auto_memory_endpoint_identity_out_3_a_bits_source,
  output [33:0]  auto_memory_endpoint_identity_out_3_a_bits_address,
  output [63:0]  auto_memory_endpoint_identity_out_3_a_bits_mask,
  output         auto_memory_endpoint_identity_out_3_d_ready,
  input          auto_memory_endpoint_identity_out_3_d_valid,
  input  [3:0]   auto_memory_endpoint_identity_out_3_d_bits_source,
  input          auto_memory_endpoint_identity_out_2_a_ready,
  output         auto_memory_endpoint_identity_out_2_a_valid,
  output [2:0]   auto_memory_endpoint_identity_out_2_a_bits_size,
  output [3:0]   auto_memory_endpoint_identity_out_2_a_bits_source,
  output [33:0]  auto_memory_endpoint_identity_out_2_a_bits_address,
  output [63:0]  auto_memory_endpoint_identity_out_2_a_bits_mask,
  output         auto_memory_endpoint_identity_out_2_d_ready,
  input          auto_memory_endpoint_identity_out_2_d_valid,
  input  [3:0]   auto_memory_endpoint_identity_out_2_d_bits_source,
  input          auto_memory_endpoint_identity_out_1_a_ready,
  output         auto_memory_endpoint_identity_out_1_a_valid,
  output [2:0]   auto_memory_endpoint_identity_out_1_a_bits_size,
  output [3:0]   auto_memory_endpoint_identity_out_1_a_bits_source,
  output [33:0]  auto_memory_endpoint_identity_out_1_a_bits_address,
  output [63:0]  auto_memory_endpoint_identity_out_1_a_bits_mask,
  output         auto_memory_endpoint_identity_out_1_d_ready,
  input          auto_memory_endpoint_identity_out_1_d_valid,
  input  [3:0]   auto_memory_endpoint_identity_out_1_d_bits_source,
  input  [511:0] auto_memory_endpoint_identity_out_1_d_bits_data,
  input          auto_memory_endpoint_identity_out_0_a_ready,
  output         auto_memory_endpoint_identity_out_0_a_valid,
  output         auto_memory_endpoint_identity_out_0_a_bits_source,
  output [33:0]  auto_memory_endpoint_identity_out_0_a_bits_address,
  output [63:0]  auto_memory_endpoint_identity_out_0_a_bits_mask,
  output [511:0] auto_memory_endpoint_identity_out_0_a_bits_data,
  output         auto_memory_endpoint_identity_out_0_d_ready,
  input          auto_memory_endpoint_identity_out_0_d_valid,
  input          auto_memory_endpoint_identity_out_0_d_bits_source,
  output         sw_io_cmd_ready,
  input          sw_io_cmd_valid,
  input  [4:0]   sw_io_cmd_bits_inst_rs1,
  input  [4:0]   sw_io_cmd_bits_inst_rs2,
  input  [2:0]   sw_io_cmd_bits_inst_funct,
  input  [7:0]   sw_io_cmd_bits_core_id,
  input  [55:0]  sw_io_cmd_bits_payload1,
  input  [63:0]  sw_io_cmd_bits_payload2,
  input          sw_io_resp_ready,
  output         sw_io_resp_valid,
  output [4:0]   sw_io_resp_bits_rd,
  output [3:0]   sw_io_resp_bits_system_id,
  output [7:0]   sw_io_resp_bits_core_id,
  output [46:0]  sw_io_resp_bits_data
);
  wire  cores_clock; // @[ComposerSystem.scala 22:15]
  wire  cores_reset; // @[ComposerSystem.scala 22:15]
  wire  cores_auto_solvated_mem_out_a_ready; // @[ComposerSystem.scala 22:15]
  wire  cores_auto_solvated_mem_out_a_valid; // @[ComposerSystem.scala 22:15]
  wire [2:0] cores_auto_solvated_mem_out_a_bits_size; // @[ComposerSystem.scala 22:15]
  wire [3:0] cores_auto_solvated_mem_out_a_bits_source; // @[ComposerSystem.scala 22:15]
  wire [33:0] cores_auto_solvated_mem_out_a_bits_address; // @[ComposerSystem.scala 22:15]
  wire [63:0] cores_auto_solvated_mem_out_a_bits_mask; // @[ComposerSystem.scala 22:15]
  wire  cores_auto_solvated_mem_out_d_ready; // @[ComposerSystem.scala 22:15]
  wire  cores_auto_solvated_mem_out_d_valid; // @[ComposerSystem.scala 22:15]
  wire [3:0] cores_auto_solvated_mem_out_d_bits_source; // @[ComposerSystem.scala 22:15]
  wire  cores_auto_nonBonded_mem_out_a_ready; // @[ComposerSystem.scala 22:15]
  wire  cores_auto_nonBonded_mem_out_a_valid; // @[ComposerSystem.scala 22:15]
  wire [2:0] cores_auto_nonBonded_mem_out_a_bits_size; // @[ComposerSystem.scala 22:15]
  wire [3:0] cores_auto_nonBonded_mem_out_a_bits_source; // @[ComposerSystem.scala 22:15]
  wire [33:0] cores_auto_nonBonded_mem_out_a_bits_address; // @[ComposerSystem.scala 22:15]
  wire [63:0] cores_auto_nonBonded_mem_out_a_bits_mask; // @[ComposerSystem.scala 22:15]
  wire  cores_auto_nonBonded_mem_out_d_ready; // @[ComposerSystem.scala 22:15]
  wire  cores_auto_nonBonded_mem_out_d_valid; // @[ComposerSystem.scala 22:15]
  wire [3:0] cores_auto_nonBonded_mem_out_d_bits_source; // @[ComposerSystem.scala 22:15]
  wire  cores_auto_halfNonBonded_mem_out_a_ready; // @[ComposerSystem.scala 22:15]
  wire  cores_auto_halfNonBonded_mem_out_a_valid; // @[ComposerSystem.scala 22:15]
  wire [2:0] cores_auto_halfNonBonded_mem_out_a_bits_size; // @[ComposerSystem.scala 22:15]
  wire [3:0] cores_auto_halfNonBonded_mem_out_a_bits_source; // @[ComposerSystem.scala 22:15]
  wire [33:0] cores_auto_halfNonBonded_mem_out_a_bits_address; // @[ComposerSystem.scala 22:15]
  wire [63:0] cores_auto_halfNonBonded_mem_out_a_bits_mask; // @[ComposerSystem.scala 22:15]
  wire  cores_auto_halfNonBonded_mem_out_d_ready; // @[ComposerSystem.scala 22:15]
  wire  cores_auto_halfNonBonded_mem_out_d_valid; // @[ComposerSystem.scala 22:15]
  wire [3:0] cores_auto_halfNonBonded_mem_out_d_bits_source; // @[ComposerSystem.scala 22:15]
  wire  cores_auto_data_mem_out_a_ready; // @[ComposerSystem.scala 22:15]
  wire  cores_auto_data_mem_out_a_valid; // @[ComposerSystem.scala 22:15]
  wire [2:0] cores_auto_data_mem_out_a_bits_size; // @[ComposerSystem.scala 22:15]
  wire [3:0] cores_auto_data_mem_out_a_bits_source; // @[ComposerSystem.scala 22:15]
  wire [33:0] cores_auto_data_mem_out_a_bits_address; // @[ComposerSystem.scala 22:15]
  wire [63:0] cores_auto_data_mem_out_a_bits_mask; // @[ComposerSystem.scala 22:15]
  wire  cores_auto_data_mem_out_d_ready; // @[ComposerSystem.scala 22:15]
  wire  cores_auto_data_mem_out_d_valid; // @[ComposerSystem.scala 22:15]
  wire [3:0] cores_auto_data_mem_out_d_bits_source; // @[ComposerSystem.scala 22:15]
  wire [511:0] cores_auto_data_mem_out_d_bits_data; // @[ComposerSystem.scala 22:15]
  wire  cores_auto_writers_out_a_ready; // @[ComposerSystem.scala 22:15]
  wire  cores_auto_writers_out_a_valid; // @[ComposerSystem.scala 22:15]
  wire  cores_auto_writers_out_a_bits_source; // @[ComposerSystem.scala 22:15]
  wire [33:0] cores_auto_writers_out_a_bits_address; // @[ComposerSystem.scala 22:15]
  wire [63:0] cores_auto_writers_out_a_bits_mask; // @[ComposerSystem.scala 22:15]
  wire [511:0] cores_auto_writers_out_a_bits_data; // @[ComposerSystem.scala 22:15]
  wire  cores_auto_writers_out_d_ready; // @[ComposerSystem.scala 22:15]
  wire  cores_auto_writers_out_d_valid; // @[ComposerSystem.scala 22:15]
  wire  cores_auto_writers_out_d_bits_source; // @[ComposerSystem.scala 22:15]
  wire  cores_io_req_ready; // @[ComposerSystem.scala 22:15]
  wire  cores_io_req_valid; // @[ComposerSystem.scala 22:15]
  wire [4:0] cores_io_req_bits_inst_rs1; // @[ComposerSystem.scala 22:15]
  wire [55:0] cores_io_req_bits_payload1; // @[ComposerSystem.scala 22:15]
  wire [63:0] cores_io_req_bits_payload2; // @[ComposerSystem.scala 22:15]
  wire  cores_io_resp_ready; // @[ComposerSystem.scala 22:15]
  wire  cores_io_resp_valid; // @[ComposerSystem.scala 22:15]
  wire  cores_myWriters_WriteChannel_valid; // @[ComposerSystem.scala 22:15]
  wire [33:0] cores_myWriters_WriteChannel_bits_addr; // @[ComposerSystem.scala 22:15]
  wire [33:0] cores_myWriters_WriteChannel_bits_len; // @[ComposerSystem.scala 22:15]
  wire  respArbiter_io_in_0_ready; // @[ComposerSystem.scala 133:27]
  wire  respArbiter_io_in_0_valid; // @[ComposerSystem.scala 133:27]
  wire [59:0] respArbiter_io_in_0_bits_data; // @[ComposerSystem.scala 133:27]
  wire [4:0] respArbiter_io_in_0_bits_rd; // @[ComposerSystem.scala 133:27]
  wire  respArbiter_io_out_ready; // @[ComposerSystem.scala 133:27]
  wire  respArbiter_io_out_valid; // @[ComposerSystem.scala 133:27]
  wire [59:0] respArbiter_io_out_bits_data; // @[ComposerSystem.scala 133:27]
  wire [4:0] respArbiter_io_out_bits_rd; // @[ComposerSystem.scala 133:27]
  wire  cmdArbiter_io_in_0_ready; // @[ComposerSystem.scala 140:26]
  wire  cmdArbiter_io_in_0_valid; // @[ComposerSystem.scala 140:26]
  wire [4:0] cmdArbiter_io_in_0_bits_inst_rs1; // @[ComposerSystem.scala 140:26]
  wire [4:0] cmdArbiter_io_in_0_bits_inst_rs2; // @[ComposerSystem.scala 140:26]
  wire [2:0] cmdArbiter_io_in_0_bits_inst_funct; // @[ComposerSystem.scala 140:26]
  wire [7:0] cmdArbiter_io_in_0_bits_core_id; // @[ComposerSystem.scala 140:26]
  wire [55:0] cmdArbiter_io_in_0_bits_payload1; // @[ComposerSystem.scala 140:26]
  wire [63:0] cmdArbiter_io_in_0_bits_payload2; // @[ComposerSystem.scala 140:26]
  wire  cmdArbiter_io_out_ready; // @[ComposerSystem.scala 140:26]
  wire  cmdArbiter_io_out_valid; // @[ComposerSystem.scala 140:26]
  wire [4:0] cmdArbiter_io_out_bits_inst_rs1; // @[ComposerSystem.scala 140:26]
  wire [4:0] cmdArbiter_io_out_bits_inst_rs2; // @[ComposerSystem.scala 140:26]
  wire [2:0] cmdArbiter_io_out_bits_inst_funct; // @[ComposerSystem.scala 140:26]
  wire [7:0] cmdArbiter_io_out_bits_core_id; // @[ComposerSystem.scala 140:26]
  wire [55:0] cmdArbiter_io_out_bits_payload1; // @[ComposerSystem.scala 140:26]
  wire [63:0] cmdArbiter_io_out_bits_payload2; // @[ComposerSystem.scala 140:26]
  wire  cmd_clock; // @[Decoupled.scala 375:21]
  wire  cmd_reset; // @[Decoupled.scala 375:21]
  wire  cmd_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  cmd_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [4:0] cmd_io_enq_bits_inst_rs1; // @[Decoupled.scala 375:21]
  wire [4:0] cmd_io_enq_bits_inst_rs2; // @[Decoupled.scala 375:21]
  wire [2:0] cmd_io_enq_bits_inst_funct; // @[Decoupled.scala 375:21]
  wire [7:0] cmd_io_enq_bits_core_id; // @[Decoupled.scala 375:21]
  wire [55:0] cmd_io_enq_bits_payload1; // @[Decoupled.scala 375:21]
  wire [63:0] cmd_io_enq_bits_payload2; // @[Decoupled.scala 375:21]
  wire  cmd_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  cmd_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [4:0] cmd_io_deq_bits_inst_rs1; // @[Decoupled.scala 375:21]
  wire [4:0] cmd_io_deq_bits_inst_rs2; // @[Decoupled.scala 375:21]
  wire [2:0] cmd_io_deq_bits_inst_funct; // @[Decoupled.scala 375:21]
  wire [7:0] cmd_io_deq_bits_core_id; // @[Decoupled.scala 375:21]
  wire [55:0] cmd_io_deq_bits_payload1; // @[Decoupled.scala 375:21]
  wire [63:0] cmd_io_deq_bits_payload2; // @[Decoupled.scala 375:21]
  wire  coreResps_rq_clock; // @[ComposerSystem.scala 212:22]
  wire  coreResps_rq_reset; // @[ComposerSystem.scala 212:22]
  wire  coreResps_rq_io_enq_ready; // @[ComposerSystem.scala 212:22]
  wire  coreResps_rq_io_enq_valid; // @[ComposerSystem.scala 212:22]
  wire  coreResps_rq_io_deq_ready; // @[ComposerSystem.scala 212:22]
  wire  coreResps_rq_io_deq_valid; // @[ComposerSystem.scala 212:22]
  wire [59:0] coreResps_rq_io_deq_bits_data; // @[ComposerSystem.scala 212:22]
  wire [4:0] coreResps_rq_io_deq_bits_rd; // @[ComposerSystem.scala 212:22]
  wire  respQ_clock; // @[Decoupled.scala 375:21]
  wire  respQ_reset; // @[Decoupled.scala 375:21]
  wire  respQ_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  respQ_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [4:0] respQ_io_enq_bits_rd; // @[Decoupled.scala 375:21]
  wire [46:0] respQ_io_enq_bits_data; // @[Decoupled.scala 375:21]
  wire  respQ_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  respQ_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [4:0] respQ_io_deq_bits_rd; // @[Decoupled.scala 375:21]
  wire [3:0] respQ_io_deq_bits_system_id; // @[Decoupled.scala 375:21]
  wire [7:0] respQ_io_deq_bits_core_id; // @[Decoupled.scala 375:21]
  wire [46:0] respQ_io_deq_bits_data; // @[Decoupled.scala 375:21]
  wire [7:0] channelSelect = {cmd_io_deq_bits_inst_rs2[2:0],cmd_io_deq_bits_inst_rs1}; // @[Cat.scala 33:92]
  wire  _coreStart_T = cmd_io_deq_ready & cmd_io_deq_valid; // @[Decoupled.scala 51:35]
  wire  _coreStart_T_3 = cmd_io_deq_bits_core_id == 8'h0; // @[ComposerSystem.scala 304:78]
  reg  cmdPipePipe_valid; // @[Valid.scala 130:22]
  reg  cmdPipePipe_bits_start; // @[Reg.scala 19:16]
  reg [4:0] cmdPipePipe_bits_cmdP_inst_rs1; // @[Reg.scala 19:16]
  reg [55:0] cmdPipePipe_bits_cmdP_payload1; // @[Reg.scala 19:16]
  reg [63:0] cmdPipePipe_bits_cmdP_payload2; // @[Reg.scala 19:16]
  reg  cmdPipePipe_valid_1; // @[Valid.scala 130:22]
  reg  cmdPipePipe_bits_1_start; // @[Reg.scala 19:16]
  reg [4:0] cmdPipePipe_bits_1_cmdP_inst_rs1; // @[Reg.scala 19:16]
  reg [55:0] cmdPipePipe_bits_1_cmdP_payload1; // @[Reg.scala 19:16]
  reg [63:0] cmdPipePipe_bits_1_cmdP_payload2; // @[Reg.scala 19:16]
  reg  cmdPipePipe_valid_2; // @[Valid.scala 130:22]
  reg  cmdPipePipe_bits_2_start; // @[Reg.scala 19:16]
  reg [4:0] cmdPipePipe_bits_2_cmdP_inst_rs1; // @[Reg.scala 19:16]
  reg [55:0] cmdPipePipe_bits_2_cmdP_payload1; // @[Reg.scala 19:16]
  reg [63:0] cmdPipePipe_bits_2_cmdP_payload2; // @[Reg.scala 19:16]
  reg  cmdPipePipe_valid_3; // @[Valid.scala 130:22]
  reg  cmdPipePipe_bits_3_start; // @[Reg.scala 19:16]
  reg [4:0] cmdPipePipe_bits_3_cmdP_inst_rs1; // @[Reg.scala 19:16]
  reg [55:0] cmdPipePipe_bits_3_cmdP_payload1; // @[Reg.scala 19:16]
  reg [63:0] cmdPipePipe_bits_3_cmdP_payload2; // @[Reg.scala 19:16]
  reg  cmdFireLatch; // @[ComposerSystem.scala 322:29]
  reg [2:0] cmdBitsLatch_inst_funct; // @[ComposerSystem.scala 323:29]
  reg [7:0] cmdBitsLatch_core_id; // @[ComposerSystem.scala 323:29]
  wire  addr_func_live = cmd_io_deq_bits_inst_funct == 3'h0 & _coreStart_T; // @[ComposerSystem.scala 327:68]
  wire [33:0] txLenFromCmd = cmd_io_deq_bits_payload1[33:0]; // @[ComposerSystem.scala 333:39]
  reg [33:0] tx_len; // @[ComposerSystem.scala 342:25]
  reg [33:0] tx_addr_start; // @[ComposerSystem.scala 343:32]
  ComposerCoreWrapper cores ( // @[ComposerSystem.scala 22:15]
    .clock(cores_clock),
    .reset(cores_reset),
    .auto_solvated_mem_out_a_ready(cores_auto_solvated_mem_out_a_ready),
    .auto_solvated_mem_out_a_valid(cores_auto_solvated_mem_out_a_valid),
    .auto_solvated_mem_out_a_bits_size(cores_auto_solvated_mem_out_a_bits_size),
    .auto_solvated_mem_out_a_bits_source(cores_auto_solvated_mem_out_a_bits_source),
    .auto_solvated_mem_out_a_bits_address(cores_auto_solvated_mem_out_a_bits_address),
    .auto_solvated_mem_out_a_bits_mask(cores_auto_solvated_mem_out_a_bits_mask),
    .auto_solvated_mem_out_d_ready(cores_auto_solvated_mem_out_d_ready),
    .auto_solvated_mem_out_d_valid(cores_auto_solvated_mem_out_d_valid),
    .auto_solvated_mem_out_d_bits_source(cores_auto_solvated_mem_out_d_bits_source),
    .auto_nonBonded_mem_out_a_ready(cores_auto_nonBonded_mem_out_a_ready),
    .auto_nonBonded_mem_out_a_valid(cores_auto_nonBonded_mem_out_a_valid),
    .auto_nonBonded_mem_out_a_bits_size(cores_auto_nonBonded_mem_out_a_bits_size),
    .auto_nonBonded_mem_out_a_bits_source(cores_auto_nonBonded_mem_out_a_bits_source),
    .auto_nonBonded_mem_out_a_bits_address(cores_auto_nonBonded_mem_out_a_bits_address),
    .auto_nonBonded_mem_out_a_bits_mask(cores_auto_nonBonded_mem_out_a_bits_mask),
    .auto_nonBonded_mem_out_d_ready(cores_auto_nonBonded_mem_out_d_ready),
    .auto_nonBonded_mem_out_d_valid(cores_auto_nonBonded_mem_out_d_valid),
    .auto_nonBonded_mem_out_d_bits_source(cores_auto_nonBonded_mem_out_d_bits_source),
    .auto_halfNonBonded_mem_out_a_ready(cores_auto_halfNonBonded_mem_out_a_ready),
    .auto_halfNonBonded_mem_out_a_valid(cores_auto_halfNonBonded_mem_out_a_valid),
    .auto_halfNonBonded_mem_out_a_bits_size(cores_auto_halfNonBonded_mem_out_a_bits_size),
    .auto_halfNonBonded_mem_out_a_bits_source(cores_auto_halfNonBonded_mem_out_a_bits_source),
    .auto_halfNonBonded_mem_out_a_bits_address(cores_auto_halfNonBonded_mem_out_a_bits_address),
    .auto_halfNonBonded_mem_out_a_bits_mask(cores_auto_halfNonBonded_mem_out_a_bits_mask),
    .auto_halfNonBonded_mem_out_d_ready(cores_auto_halfNonBonded_mem_out_d_ready),
    .auto_halfNonBonded_mem_out_d_valid(cores_auto_halfNonBonded_mem_out_d_valid),
    .auto_halfNonBonded_mem_out_d_bits_source(cores_auto_halfNonBonded_mem_out_d_bits_source),
    .auto_data_mem_out_a_ready(cores_auto_data_mem_out_a_ready),
    .auto_data_mem_out_a_valid(cores_auto_data_mem_out_a_valid),
    .auto_data_mem_out_a_bits_size(cores_auto_data_mem_out_a_bits_size),
    .auto_data_mem_out_a_bits_source(cores_auto_data_mem_out_a_bits_source),
    .auto_data_mem_out_a_bits_address(cores_auto_data_mem_out_a_bits_address),
    .auto_data_mem_out_a_bits_mask(cores_auto_data_mem_out_a_bits_mask),
    .auto_data_mem_out_d_ready(cores_auto_data_mem_out_d_ready),
    .auto_data_mem_out_d_valid(cores_auto_data_mem_out_d_valid),
    .auto_data_mem_out_d_bits_source(cores_auto_data_mem_out_d_bits_source),
    .auto_data_mem_out_d_bits_data(cores_auto_data_mem_out_d_bits_data),
    .auto_writers_out_a_ready(cores_auto_writers_out_a_ready),
    .auto_writers_out_a_valid(cores_auto_writers_out_a_valid),
    .auto_writers_out_a_bits_source(cores_auto_writers_out_a_bits_source),
    .auto_writers_out_a_bits_address(cores_auto_writers_out_a_bits_address),
    .auto_writers_out_a_bits_mask(cores_auto_writers_out_a_bits_mask),
    .auto_writers_out_a_bits_data(cores_auto_writers_out_a_bits_data),
    .auto_writers_out_d_ready(cores_auto_writers_out_d_ready),
    .auto_writers_out_d_valid(cores_auto_writers_out_d_valid),
    .auto_writers_out_d_bits_source(cores_auto_writers_out_d_bits_source),
    .io_req_ready(cores_io_req_ready),
    .io_req_valid(cores_io_req_valid),
    .io_req_bits_inst_rs1(cores_io_req_bits_inst_rs1),
    .io_req_bits_payload1(cores_io_req_bits_payload1),
    .io_req_bits_payload2(cores_io_req_bits_payload2),
    .io_resp_ready(cores_io_resp_ready),
    .io_resp_valid(cores_io_resp_valid),
    .myWriters_WriteChannel_valid(cores_myWriters_WriteChannel_valid),
    .myWriters_WriteChannel_bits_addr(cores_myWriters_WriteChannel_bits_addr),
    .myWriters_WriteChannel_bits_len(cores_myWriters_WriteChannel_bits_len)
  );
  MultiLevelArbiter respArbiter ( // @[ComposerSystem.scala 133:27]
    .io_in_0_ready(respArbiter_io_in_0_ready),
    .io_in_0_valid(respArbiter_io_in_0_valid),
    .io_in_0_bits_data(respArbiter_io_in_0_bits_data),
    .io_in_0_bits_rd(respArbiter_io_in_0_bits_rd),
    .io_out_ready(respArbiter_io_out_ready),
    .io_out_valid(respArbiter_io_out_valid),
    .io_out_bits_data(respArbiter_io_out_bits_data),
    .io_out_bits_rd(respArbiter_io_out_bits_rd)
  );
  RRArbiter cmdArbiter ( // @[ComposerSystem.scala 140:26]
    .io_in_0_ready(cmdArbiter_io_in_0_ready),
    .io_in_0_valid(cmdArbiter_io_in_0_valid),
    .io_in_0_bits_inst_rs1(cmdArbiter_io_in_0_bits_inst_rs1),
    .io_in_0_bits_inst_rs2(cmdArbiter_io_in_0_bits_inst_rs2),
    .io_in_0_bits_inst_funct(cmdArbiter_io_in_0_bits_inst_funct),
    .io_in_0_bits_core_id(cmdArbiter_io_in_0_bits_core_id),
    .io_in_0_bits_payload1(cmdArbiter_io_in_0_bits_payload1),
    .io_in_0_bits_payload2(cmdArbiter_io_in_0_bits_payload2),
    .io_out_ready(cmdArbiter_io_out_ready),
    .io_out_valid(cmdArbiter_io_out_valid),
    .io_out_bits_inst_rs1(cmdArbiter_io_out_bits_inst_rs1),
    .io_out_bits_inst_rs2(cmdArbiter_io_out_bits_inst_rs2),
    .io_out_bits_inst_funct(cmdArbiter_io_out_bits_inst_funct),
    .io_out_bits_core_id(cmdArbiter_io_out_bits_core_id),
    .io_out_bits_payload1(cmdArbiter_io_out_bits_payload1),
    .io_out_bits_payload2(cmdArbiter_io_out_bits_payload2)
  );
  Queue cmd ( // @[Decoupled.scala 375:21]
    .clock(cmd_clock),
    .reset(cmd_reset),
    .io_enq_ready(cmd_io_enq_ready),
    .io_enq_valid(cmd_io_enq_valid),
    .io_enq_bits_inst_rs1(cmd_io_enq_bits_inst_rs1),
    .io_enq_bits_inst_rs2(cmd_io_enq_bits_inst_rs2),
    .io_enq_bits_inst_funct(cmd_io_enq_bits_inst_funct),
    .io_enq_bits_core_id(cmd_io_enq_bits_core_id),
    .io_enq_bits_payload1(cmd_io_enq_bits_payload1),
    .io_enq_bits_payload2(cmd_io_enq_bits_payload2),
    .io_deq_ready(cmd_io_deq_ready),
    .io_deq_valid(cmd_io_deq_valid),
    .io_deq_bits_inst_rs1(cmd_io_deq_bits_inst_rs1),
    .io_deq_bits_inst_rs2(cmd_io_deq_bits_inst_rs2),
    .io_deq_bits_inst_funct(cmd_io_deq_bits_inst_funct),
    .io_deq_bits_core_id(cmd_io_deq_bits_core_id),
    .io_deq_bits_payload1(cmd_io_deq_bits_payload1),
    .io_deq_bits_payload2(cmd_io_deq_bits_payload2)
  );
  Queue_1 coreResps_rq ( // @[ComposerSystem.scala 212:22]
    .clock(coreResps_rq_clock),
    .reset(coreResps_rq_reset),
    .io_enq_ready(coreResps_rq_io_enq_ready),
    .io_enq_valid(coreResps_rq_io_enq_valid),
    .io_deq_ready(coreResps_rq_io_deq_ready),
    .io_deq_valid(coreResps_rq_io_deq_valid),
    .io_deq_bits_data(coreResps_rq_io_deq_bits_data),
    .io_deq_bits_rd(coreResps_rq_io_deq_bits_rd)
  );
  Queue_2 respQ ( // @[Decoupled.scala 375:21]
    .clock(respQ_clock),
    .reset(respQ_reset),
    .io_enq_ready(respQ_io_enq_ready),
    .io_enq_valid(respQ_io_enq_valid),
    .io_enq_bits_rd(respQ_io_enq_bits_rd),
    .io_enq_bits_data(respQ_io_enq_bits_data),
    .io_deq_ready(respQ_io_deq_ready),
    .io_deq_valid(respQ_io_deq_valid),
    .io_deq_bits_rd(respQ_io_deq_bits_rd),
    .io_deq_bits_system_id(respQ_io_deq_bits_system_id),
    .io_deq_bits_core_id(respQ_io_deq_bits_core_id),
    .io_deq_bits_data(respQ_io_deq_bits_data)
  );
  assign auto_memory_endpoint_identity_out_4_a_valid = cores_auto_solvated_mem_out_a_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_4_a_bits_size = cores_auto_solvated_mem_out_a_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_4_a_bits_source = cores_auto_solvated_mem_out_a_bits_source; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_4_a_bits_address = cores_auto_solvated_mem_out_a_bits_address; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_4_a_bits_mask = cores_auto_solvated_mem_out_a_bits_mask; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_4_d_ready = cores_auto_solvated_mem_out_d_ready; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_3_a_valid = cores_auto_nonBonded_mem_out_a_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_3_a_bits_size = cores_auto_nonBonded_mem_out_a_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_3_a_bits_source = cores_auto_nonBonded_mem_out_a_bits_source; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_3_a_bits_address = cores_auto_nonBonded_mem_out_a_bits_address; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_3_a_bits_mask = cores_auto_nonBonded_mem_out_a_bits_mask; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_3_d_ready = cores_auto_nonBonded_mem_out_d_ready; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_2_a_valid = cores_auto_halfNonBonded_mem_out_a_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_2_a_bits_size = cores_auto_halfNonBonded_mem_out_a_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_2_a_bits_source = cores_auto_halfNonBonded_mem_out_a_bits_source; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_2_a_bits_address = cores_auto_halfNonBonded_mem_out_a_bits_address; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_2_a_bits_mask = cores_auto_halfNonBonded_mem_out_a_bits_mask; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_2_d_ready = cores_auto_halfNonBonded_mem_out_d_ready; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_1_a_valid = cores_auto_data_mem_out_a_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_1_a_bits_size = cores_auto_data_mem_out_a_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_1_a_bits_source = cores_auto_data_mem_out_a_bits_source; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_1_a_bits_address = cores_auto_data_mem_out_a_bits_address; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_1_a_bits_mask = cores_auto_data_mem_out_a_bits_mask; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_1_d_ready = cores_auto_data_mem_out_d_ready; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_0_a_valid = cores_auto_writers_out_a_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_0_a_bits_source = cores_auto_writers_out_a_bits_source; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_0_a_bits_address = cores_auto_writers_out_a_bits_address; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_0_a_bits_mask = cores_auto_writers_out_a_bits_mask; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_0_a_bits_data = cores_auto_writers_out_a_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_memory_endpoint_identity_out_0_d_ready = cores_auto_writers_out_d_ready; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign sw_io_cmd_ready = cmdArbiter_io_in_0_ready; // @[ComposerSystem.scala 156:21 166:27]
  assign sw_io_resp_valid = respQ_io_deq_valid; // @[ComposerSystem.scala 278:20]
  assign sw_io_resp_bits_rd = respQ_io_deq_bits_rd; // @[ComposerSystem.scala 278:20]
  assign sw_io_resp_bits_system_id = respQ_io_deq_bits_system_id; // @[ComposerSystem.scala 278:20]
  assign sw_io_resp_bits_core_id = respQ_io_deq_bits_core_id; // @[ComposerSystem.scala 278:20]
  assign sw_io_resp_bits_data = respQ_io_deq_bits_data; // @[ComposerSystem.scala 278:20]
  assign cores_clock = clock;
  assign cores_reset = reset;
  assign cores_auto_solvated_mem_out_a_ready = auto_memory_endpoint_identity_out_4_a_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign cores_auto_solvated_mem_out_d_valid = auto_memory_endpoint_identity_out_4_d_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign cores_auto_solvated_mem_out_d_bits_source = auto_memory_endpoint_identity_out_4_d_bits_source; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign cores_auto_nonBonded_mem_out_a_ready = auto_memory_endpoint_identity_out_3_a_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign cores_auto_nonBonded_mem_out_d_valid = auto_memory_endpoint_identity_out_3_d_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign cores_auto_nonBonded_mem_out_d_bits_source = auto_memory_endpoint_identity_out_3_d_bits_source; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign cores_auto_halfNonBonded_mem_out_a_ready = auto_memory_endpoint_identity_out_2_a_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign cores_auto_halfNonBonded_mem_out_d_valid = auto_memory_endpoint_identity_out_2_d_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign cores_auto_halfNonBonded_mem_out_d_bits_source = auto_memory_endpoint_identity_out_2_d_bits_source; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign cores_auto_data_mem_out_a_ready = auto_memory_endpoint_identity_out_1_a_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign cores_auto_data_mem_out_d_valid = auto_memory_endpoint_identity_out_1_d_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign cores_auto_data_mem_out_d_bits_source = auto_memory_endpoint_identity_out_1_d_bits_source; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign cores_auto_data_mem_out_d_bits_data = auto_memory_endpoint_identity_out_1_d_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign cores_auto_writers_out_a_ready = auto_memory_endpoint_identity_out_0_a_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign cores_auto_writers_out_d_valid = auto_memory_endpoint_identity_out_0_d_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign cores_auto_writers_out_d_bits_source = auto_memory_endpoint_identity_out_0_d_bits_source; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign cores_io_req_valid = cmdPipePipe_bits_3_start & cmdPipePipe_valid_3; // @[ComposerSystem.scala 313:47]
  assign cores_io_req_bits_inst_rs1 = cmdPipePipe_bits_3_cmdP_inst_rs1; // @[Valid.scala 125:21 127:16]
  assign cores_io_req_bits_payload1 = cmdPipePipe_bits_3_cmdP_payload1; // @[Valid.scala 125:21 127:16]
  assign cores_io_req_bits_payload2 = cmdPipePipe_bits_3_cmdP_payload2; // @[Valid.scala 125:21 127:16]
  assign cores_io_resp_ready = coreResps_rq_io_enq_ready; // @[ComposerSystem.scala 213:17]
  assign cores_myWriters_WriteChannel_valid = cmdFireLatch & cmdBitsLatch_inst_funct == 3'h1 & cmdBitsLatch_core_id == 8'h0
    ; // @[ComposerSystem.scala 348:75]
  assign cores_myWriters_WriteChannel_bits_addr = tx_addr_start; // @[ComposerSystem.scala 349:24]
  assign cores_myWriters_WriteChannel_bits_len = tx_len; // @[ComposerSystem.scala 350:23]
  assign respArbiter_io_in_0_valid = coreResps_rq_io_deq_valid; // @[ComposerSystem.scala 219:21]
  assign respArbiter_io_in_0_bits_data = coreResps_rq_io_deq_bits_data; // @[ComposerSystem.scala 219:21]
  assign respArbiter_io_in_0_bits_rd = coreResps_rq_io_deq_bits_rd; // @[ComposerSystem.scala 219:21]
  assign respArbiter_io_out_ready = respQ_io_enq_ready; // @[ComposerSystem.scala 220:18 Decoupled.scala 379:17]
  assign cmdArbiter_io_in_0_valid = sw_io_cmd_valid; // @[ComposerSystem.scala 156:21 158:17]
  assign cmdArbiter_io_in_0_bits_inst_rs1 = sw_io_cmd_bits_inst_rs1; // @[ComposerSystem.scala 156:21 160:16]
  assign cmdArbiter_io_in_0_bits_inst_rs2 = sw_io_cmd_bits_inst_rs2; // @[ComposerSystem.scala 156:21 160:16]
  assign cmdArbiter_io_in_0_bits_inst_funct = sw_io_cmd_bits_inst_funct; // @[ComposerSystem.scala 156:21 160:16]
  assign cmdArbiter_io_in_0_bits_core_id = sw_io_cmd_bits_core_id; // @[ComposerSystem.scala 156:21 160:16]
  assign cmdArbiter_io_in_0_bits_payload1 = sw_io_cmd_bits_payload1; // @[ComposerSystem.scala 156:21 160:16]
  assign cmdArbiter_io_in_0_bits_payload2 = sw_io_cmd_bits_payload2; // @[ComposerSystem.scala 156:21 160:16]
  assign cmdArbiter_io_out_ready = cmd_io_enq_ready; // @[Decoupled.scala 379:17]
  assign cmd_clock = clock;
  assign cmd_reset = reset;
  assign cmd_io_enq_valid = cmdArbiter_io_out_valid; // @[Decoupled.scala 377:22]
  assign cmd_io_enq_bits_inst_rs1 = cmdArbiter_io_out_bits_inst_rs1; // @[Decoupled.scala 378:21]
  assign cmd_io_enq_bits_inst_rs2 = cmdArbiter_io_out_bits_inst_rs2; // @[Decoupled.scala 378:21]
  assign cmd_io_enq_bits_inst_funct = cmdArbiter_io_out_bits_inst_funct; // @[Decoupled.scala 378:21]
  assign cmd_io_enq_bits_core_id = cmdArbiter_io_out_bits_core_id; // @[Decoupled.scala 378:21]
  assign cmd_io_enq_bits_payload1 = cmdArbiter_io_out_bits_payload1; // @[Decoupled.scala 378:21]
  assign cmd_io_enq_bits_payload2 = cmdArbiter_io_out_bits_payload2; // @[Decoupled.scala 378:21]
  assign cmd_io_deq_ready = cmd_io_deq_bits_inst_funct != 3'h1 | cores_io_req_ready; // @[ComposerSystem.scala 194:47]
  assign coreResps_rq_clock = clock;
  assign coreResps_rq_reset = reset;
  assign coreResps_rq_io_enq_valid = cores_io_resp_valid; // @[ComposerSystem.scala 213:17]
  assign coreResps_rq_io_deq_ready = respArbiter_io_in_0_ready; // @[ComposerSystem.scala 219:21]
  assign respQ_clock = clock;
  assign respQ_reset = reset;
  assign respQ_io_enq_valid = respArbiter_io_out_valid; // @[ComposerSystem.scala 220:18 221:14]
  assign respQ_io_enq_bits_rd = respArbiter_io_out_bits_rd; // @[ComposerSystem.scala 220:18 222:16]
  assign respQ_io_enq_bits_data = respArbiter_io_out_bits_data[46:0]; // @[ComposerSystem.scala 220:18 224:18]
  assign respQ_io_deq_ready = sw_io_resp_ready; // @[ComposerSystem.scala 278:20]
  always @(posedge clock) begin
    if (reset) begin // @[Valid.scala 130:22]
      cmdPipePipe_valid <= 1'h0; // @[Valid.scala 130:22]
    end else begin
      cmdPipePipe_valid <= 1'h1; // @[Valid.scala 130:22]
    end
    cmdPipePipe_bits_start <= _coreStart_T & cmd_io_deq_bits_inst_funct == 3'h1 & cmd_io_deq_bits_core_id == 8'h0; // @[ComposerSystem.scala 304:64]
    cmdPipePipe_bits_cmdP_inst_rs1 <= cmd_io_deq_bits_inst_rs1; // @[ComposerSystem.scala 306:24 312:19]
    cmdPipePipe_bits_cmdP_payload1 <= cmd_io_deq_bits_payload1; // @[ComposerSystem.scala 306:24 312:19]
    cmdPipePipe_bits_cmdP_payload2 <= cmd_io_deq_bits_payload2; // @[ComposerSystem.scala 306:24 312:19]
    if (reset) begin // @[Valid.scala 130:22]
      cmdPipePipe_valid_1 <= 1'h0; // @[Valid.scala 130:22]
    end else begin
      cmdPipePipe_valid_1 <= cmdPipePipe_valid; // @[Valid.scala 130:22]
    end
    if (cmdPipePipe_valid) begin // @[Reg.scala 20:18]
      cmdPipePipe_bits_1_start <= cmdPipePipe_bits_start; // @[Reg.scala 20:22]
    end
    if (cmdPipePipe_valid) begin // @[Reg.scala 20:18]
      cmdPipePipe_bits_1_cmdP_inst_rs1 <= cmdPipePipe_bits_cmdP_inst_rs1; // @[Reg.scala 20:22]
    end
    if (cmdPipePipe_valid) begin // @[Reg.scala 20:18]
      cmdPipePipe_bits_1_cmdP_payload1 <= cmdPipePipe_bits_cmdP_payload1; // @[Reg.scala 20:22]
    end
    if (cmdPipePipe_valid) begin // @[Reg.scala 20:18]
      cmdPipePipe_bits_1_cmdP_payload2 <= cmdPipePipe_bits_cmdP_payload2; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[Valid.scala 130:22]
      cmdPipePipe_valid_2 <= 1'h0; // @[Valid.scala 130:22]
    end else begin
      cmdPipePipe_valid_2 <= cmdPipePipe_valid_1; // @[Valid.scala 130:22]
    end
    if (cmdPipePipe_valid_1) begin // @[Reg.scala 20:18]
      cmdPipePipe_bits_2_start <= cmdPipePipe_bits_1_start; // @[Reg.scala 20:22]
    end
    if (cmdPipePipe_valid_1) begin // @[Reg.scala 20:18]
      cmdPipePipe_bits_2_cmdP_inst_rs1 <= cmdPipePipe_bits_1_cmdP_inst_rs1; // @[Reg.scala 20:22]
    end
    if (cmdPipePipe_valid_1) begin // @[Reg.scala 20:18]
      cmdPipePipe_bits_2_cmdP_payload1 <= cmdPipePipe_bits_1_cmdP_payload1; // @[Reg.scala 20:22]
    end
    if (cmdPipePipe_valid_1) begin // @[Reg.scala 20:18]
      cmdPipePipe_bits_2_cmdP_payload2 <= cmdPipePipe_bits_1_cmdP_payload2; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[Valid.scala 130:22]
      cmdPipePipe_valid_3 <= 1'h0; // @[Valid.scala 130:22]
    end else begin
      cmdPipePipe_valid_3 <= cmdPipePipe_valid_2; // @[Valid.scala 130:22]
    end
    if (cmdPipePipe_valid_2) begin // @[Reg.scala 20:18]
      cmdPipePipe_bits_3_start <= cmdPipePipe_bits_2_start; // @[Reg.scala 20:22]
    end
    if (cmdPipePipe_valid_2) begin // @[Reg.scala 20:18]
      cmdPipePipe_bits_3_cmdP_inst_rs1 <= cmdPipePipe_bits_2_cmdP_inst_rs1; // @[Reg.scala 20:22]
    end
    if (cmdPipePipe_valid_2) begin // @[Reg.scala 20:18]
      cmdPipePipe_bits_3_cmdP_payload1 <= cmdPipePipe_bits_2_cmdP_payload1; // @[Reg.scala 20:22]
    end
    if (cmdPipePipe_valid_2) begin // @[Reg.scala 20:18]
      cmdPipePipe_bits_3_cmdP_payload2 <= cmdPipePipe_bits_2_cmdP_payload2; // @[Reg.scala 20:22]
    end
    cmdFireLatch <= cmd_io_deq_ready & cmd_io_deq_valid; // @[Decoupled.scala 51:35]
    cmdBitsLatch_inst_funct <= cmd_io_deq_bits_inst_funct; // @[ComposerSystem.scala 323:29]
    cmdBitsLatch_core_id <= cmd_io_deq_bits_core_id; // @[ComposerSystem.scala 323:29]
    if (addr_func_live & _coreStart_T_3 & channelSelect == 8'h0) begin // @[ComposerSystem.scala 344:91]
      tx_len <= txLenFromCmd; // @[ComposerSystem.scala 345:18]
    end
    if (addr_func_live & _coreStart_T_3 & channelSelect == 8'h0) begin // @[ComposerSystem.scala 344:91]
      tx_addr_start <= cmd_io_deq_bits_payload2[33:0]; // @[ComposerSystem.scala 346:25]
    end
  end
endmodule
module Queue_3(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [6:0]  io_enq_bits_inst_funct,
  input  [4:0]  io_enq_bits_inst_rs2,
  input  [4:0]  io_enq_bits_inst_rs1,
  input  [6:0]  io_enq_bits_inst_opcode,
  input  [63:0] io_enq_bits_rs1,
  input  [63:0] io_enq_bits_rs2,
  input         io_deq_ready,
  output        io_deq_valid,
  output [6:0]  io_deq_bits_inst_funct,
  output [4:0]  io_deq_bits_inst_rs2,
  output [4:0]  io_deq_bits_inst_rs1,
  output [6:0]  io_deq_bits_inst_opcode,
  output [63:0] io_deq_bits_rs1,
  output [63:0] io_deq_bits_rs2
);
  reg [6:0] ram_inst_funct [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_inst_funct_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_inst_funct_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [6:0] ram_inst_funct_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [6:0] ram_inst_funct_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_inst_funct_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_inst_funct_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_inst_funct_MPORT_en; // @[Decoupled.scala 273:95]
  reg [4:0] ram_inst_rs2 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_inst_rs2_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_inst_rs2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [4:0] ram_inst_rs2_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [4:0] ram_inst_rs2_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_inst_rs2_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_inst_rs2_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_inst_rs2_MPORT_en; // @[Decoupled.scala 273:95]
  reg [4:0] ram_inst_rs1 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_inst_rs1_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_inst_rs1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [4:0] ram_inst_rs1_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [4:0] ram_inst_rs1_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_inst_rs1_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_inst_rs1_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_inst_rs1_MPORT_en; // @[Decoupled.scala 273:95]
  reg [6:0] ram_inst_opcode [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_inst_opcode_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_inst_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [6:0] ram_inst_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [6:0] ram_inst_opcode_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_inst_opcode_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_inst_opcode_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_inst_opcode_MPORT_en; // @[Decoupled.scala 273:95]
  reg [63:0] ram_rs1 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_rs1_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_rs1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [63:0] ram_rs1_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [63:0] ram_rs1_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_rs1_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_rs1_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_rs1_MPORT_en; // @[Decoupled.scala 273:95]
  reg [63:0] ram_rs2 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_rs2_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_rs2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [63:0] ram_rs2_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [63:0] ram_rs2_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_rs2_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_rs2_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_rs2_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_inst_funct_io_deq_bits_MPORT_en = 1'h1;
  assign ram_inst_funct_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_inst_funct_io_deq_bits_MPORT_data = ram_inst_funct[ram_inst_funct_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_inst_funct_MPORT_data = io_enq_bits_inst_funct;
  assign ram_inst_funct_MPORT_addr = enq_ptr_value;
  assign ram_inst_funct_MPORT_mask = 1'h1;
  assign ram_inst_funct_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_inst_rs2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_inst_rs2_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_inst_rs2_io_deq_bits_MPORT_data = ram_inst_rs2[ram_inst_rs2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_inst_rs2_MPORT_data = io_enq_bits_inst_rs2;
  assign ram_inst_rs2_MPORT_addr = enq_ptr_value;
  assign ram_inst_rs2_MPORT_mask = 1'h1;
  assign ram_inst_rs2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_inst_rs1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_inst_rs1_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_inst_rs1_io_deq_bits_MPORT_data = ram_inst_rs1[ram_inst_rs1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_inst_rs1_MPORT_data = io_enq_bits_inst_rs1;
  assign ram_inst_rs1_MPORT_addr = enq_ptr_value;
  assign ram_inst_rs1_MPORT_mask = 1'h1;
  assign ram_inst_rs1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_inst_opcode_io_deq_bits_MPORT_en = 1'h1;
  assign ram_inst_opcode_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_inst_opcode_io_deq_bits_MPORT_data = ram_inst_opcode[ram_inst_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_inst_opcode_MPORT_data = io_enq_bits_inst_opcode;
  assign ram_inst_opcode_MPORT_addr = enq_ptr_value;
  assign ram_inst_opcode_MPORT_mask = 1'h1;
  assign ram_inst_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_rs1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_rs1_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_rs1_io_deq_bits_MPORT_data = ram_rs1[ram_rs1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_rs1_MPORT_data = io_enq_bits_rs1;
  assign ram_rs1_MPORT_addr = enq_ptr_value;
  assign ram_rs1_MPORT_mask = 1'h1;
  assign ram_rs1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_rs2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_rs2_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_rs2_io_deq_bits_MPORT_data = ram_rs2[ram_rs2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_rs2_MPORT_data = io_enq_bits_rs2;
  assign ram_rs2_MPORT_addr = enq_ptr_value;
  assign ram_rs2_MPORT_mask = 1'h1;
  assign ram_rs2_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_inst_funct = ram_inst_funct_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_inst_rs2 = ram_inst_rs2_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_inst_rs1 = ram_inst_rs1_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_inst_opcode = ram_inst_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_rs1 = ram_rs1_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_rs2 = ram_rs2_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_inst_funct_MPORT_en & ram_inst_funct_MPORT_mask) begin
      ram_inst_funct[ram_inst_funct_MPORT_addr] <= ram_inst_funct_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_inst_rs2_MPORT_en & ram_inst_rs2_MPORT_mask) begin
      ram_inst_rs2[ram_inst_rs2_MPORT_addr] <= ram_inst_rs2_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_inst_rs1_MPORT_en & ram_inst_rs1_MPORT_mask) begin
      ram_inst_rs1[ram_inst_rs1_MPORT_addr] <= ram_inst_rs1_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_inst_opcode_MPORT_en & ram_inst_opcode_MPORT_mask) begin
      ram_inst_opcode[ram_inst_opcode_MPORT_addr] <= ram_inst_opcode_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_rs1_MPORT_en & ram_rs1_MPORT_mask) begin
      ram_rs1[ram_rs1_MPORT_addr] <= ram_rs1_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_rs2_MPORT_en & ram_rs2_MPORT_mask) begin
      ram_rs2[ram_rs2_MPORT_addr] <= ram_rs2_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
endmodule
module RRArbiter_1(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [6:0]  io_in_0_bits_inst_funct,
  input  [4:0]  io_in_0_bits_inst_rs2,
  input  [4:0]  io_in_0_bits_inst_rs1,
  input  [6:0]  io_in_0_bits_inst_opcode,
  input  [63:0] io_in_0_bits_rs1,
  input  [63:0] io_in_0_bits_rs2,
  input         io_out_ready,
  output        io_out_valid,
  output [6:0]  io_out_bits_inst_funct,
  output [4:0]  io_out_bits_inst_rs2,
  output [4:0]  io_out_bits_inst_rs1,
  output [6:0]  io_out_bits_inst_opcode,
  output [63:0] io_out_bits_rs1,
  output [63:0] io_out_bits_rs2
);
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 74:21]
  assign io_out_valid = io_in_0_valid; // @[Arbiter.scala 55:16]
  assign io_out_bits_inst_funct = io_in_0_bits_inst_funct; // @[Arbiter.scala 56:15]
  assign io_out_bits_inst_rs2 = io_in_0_bits_inst_rs2; // @[Arbiter.scala 56:15]
  assign io_out_bits_inst_rs1 = io_in_0_bits_inst_rs1; // @[Arbiter.scala 56:15]
  assign io_out_bits_inst_opcode = io_in_0_bits_inst_opcode; // @[Arbiter.scala 56:15]
  assign io_out_bits_rs1 = io_in_0_bits_rs1; // @[Arbiter.scala 56:15]
  assign io_out_bits_rs2 = io_in_0_bits_rs2; // @[Arbiter.scala 56:15]
endmodule
module RoccCommandRouter(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [6:0]  io_in_bits_inst_funct,
  input  [4:0]  io_in_bits_inst_rs2,
  input  [4:0]  io_in_bits_inst_rs1,
  input  [6:0]  io_in_bits_inst_opcode,
  input  [63:0] io_in_bits_rs1,
  input  [63:0] io_in_bits_rs2,
  input         io_out_0_ready,
  output        io_out_0_valid,
  input         io_out_1_ready,
  output        io_out_1_valid,
  output [6:0]  io_out_1_bits_inst_funct,
  output [4:0]  io_out_1_bits_inst_rs2,
  output [4:0]  io_out_1_bits_inst_rs1,
  output [63:0] io_out_1_bits_rs1,
  output [63:0] io_out_1_bits_rs2
);
  wire  cmd_clock; // @[Decoupled.scala 375:21]
  wire  cmd_reset; // @[Decoupled.scala 375:21]
  wire  cmd_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  cmd_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [6:0] cmd_io_enq_bits_inst_funct; // @[Decoupled.scala 375:21]
  wire [4:0] cmd_io_enq_bits_inst_rs2; // @[Decoupled.scala 375:21]
  wire [4:0] cmd_io_enq_bits_inst_rs1; // @[Decoupled.scala 375:21]
  wire [6:0] cmd_io_enq_bits_inst_opcode; // @[Decoupled.scala 375:21]
  wire [63:0] cmd_io_enq_bits_rs1; // @[Decoupled.scala 375:21]
  wire [63:0] cmd_io_enq_bits_rs2; // @[Decoupled.scala 375:21]
  wire  cmd_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  cmd_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [6:0] cmd_io_deq_bits_inst_funct; // @[Decoupled.scala 375:21]
  wire [4:0] cmd_io_deq_bits_inst_rs2; // @[Decoupled.scala 375:21]
  wire [4:0] cmd_io_deq_bits_inst_rs1; // @[Decoupled.scala 375:21]
  wire [6:0] cmd_io_deq_bits_inst_opcode; // @[Decoupled.scala 375:21]
  wire [63:0] cmd_io_deq_bits_rs1; // @[Decoupled.scala 375:21]
  wire [63:0] cmd_io_deq_bits_rs2; // @[Decoupled.scala 375:21]
  wire  cmdReadys_me = 7'hb == cmd_io_deq_bits_inst_opcode; // @[LazyRoCC.scala 390:41]
  wire  cmdReadys_0 = io_out_0_ready & cmdReadys_me; // @[LazyRoCC.scala 414:15]
  wire  cmdReadys_me_1 = 7'h7b == cmd_io_deq_bits_inst_opcode; // @[LazyRoCC.scala 390:41]
  wire  cmdReadys_1 = io_out_1_ready & cmdReadys_me_1; // @[LazyRoCC.scala 414:15]
  wire [1:0] _T = cmdReadys_0 + cmdReadys_1; // @[Bitwise.scala 51:90]
  Queue_3 cmd ( // @[Decoupled.scala 375:21]
    .clock(cmd_clock),
    .reset(cmd_reset),
    .io_enq_ready(cmd_io_enq_ready),
    .io_enq_valid(cmd_io_enq_valid),
    .io_enq_bits_inst_funct(cmd_io_enq_bits_inst_funct),
    .io_enq_bits_inst_rs2(cmd_io_enq_bits_inst_rs2),
    .io_enq_bits_inst_rs1(cmd_io_enq_bits_inst_rs1),
    .io_enq_bits_inst_opcode(cmd_io_enq_bits_inst_opcode),
    .io_enq_bits_rs1(cmd_io_enq_bits_rs1),
    .io_enq_bits_rs2(cmd_io_enq_bits_rs2),
    .io_deq_ready(cmd_io_deq_ready),
    .io_deq_valid(cmd_io_deq_valid),
    .io_deq_bits_inst_funct(cmd_io_deq_bits_inst_funct),
    .io_deq_bits_inst_rs2(cmd_io_deq_bits_inst_rs2),
    .io_deq_bits_inst_rs1(cmd_io_deq_bits_inst_rs1),
    .io_deq_bits_inst_opcode(cmd_io_deq_bits_inst_opcode),
    .io_deq_bits_rs1(cmd_io_deq_bits_rs1),
    .io_deq_bits_rs2(cmd_io_deq_bits_rs2)
  );
  assign io_in_ready = cmd_io_enq_ready; // @[Decoupled.scala 379:17]
  assign io_out_0_valid = cmd_io_deq_valid & cmdReadys_me; // @[LazyRoCC.scala 412:28]
  assign io_out_1_valid = cmd_io_deq_valid & cmdReadys_me_1; // @[LazyRoCC.scala 412:28]
  assign io_out_1_bits_inst_funct = cmd_io_deq_bits_inst_funct; // @[LazyRoCC.scala 413:14]
  assign io_out_1_bits_inst_rs2 = cmd_io_deq_bits_inst_rs2; // @[LazyRoCC.scala 413:14]
  assign io_out_1_bits_inst_rs1 = cmd_io_deq_bits_inst_rs1; // @[LazyRoCC.scala 413:14]
  assign io_out_1_bits_rs1 = cmd_io_deq_bits_rs1; // @[LazyRoCC.scala 413:14]
  assign io_out_1_bits_rs2 = cmd_io_deq_bits_rs2; // @[LazyRoCC.scala 413:14]
  assign cmd_clock = clock;
  assign cmd_reset = reset;
  assign cmd_io_enq_valid = io_in_valid; // @[Decoupled.scala 377:22]
  assign cmd_io_enq_bits_inst_funct = io_in_bits_inst_funct; // @[Decoupled.scala 378:21]
  assign cmd_io_enq_bits_inst_rs2 = io_in_bits_inst_rs2; // @[Decoupled.scala 378:21]
  assign cmd_io_enq_bits_inst_rs1 = io_in_bits_inst_rs1; // @[Decoupled.scala 378:21]
  assign cmd_io_enq_bits_inst_opcode = io_in_bits_inst_opcode; // @[Decoupled.scala 378:21]
  assign cmd_io_enq_bits_rs1 = io_in_bits_rs1; // @[Decoupled.scala 378:21]
  assign cmd_io_enq_bits_rs2 = io_in_bits_rs2; // @[Decoupled.scala 378:21]
  assign cmd_io_deq_ready = cmdReadys_0 | cmdReadys_1; // @[LazyRoCC.scala 416:35]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(_T <= 2'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Custom opcode matched for more than one accelerator\n    at LazyRoCC.scala:419 assert(PopCount(cmdReadys) <= 1.U,\n"
            ); // @[LazyRoCC.scala 419:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T <= 2'h1) & ~reset) begin
          $fatal; // @[LazyRoCC.scala 419:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module RRArbiter_2(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [4:0]  io_in_0_bits_rd,
  input  [63:0] io_in_0_bits_data,
  input         io_out_ready,
  output        io_out_valid,
  output [4:0]  io_out_bits_rd,
  output [63:0] io_out_bits_data
);
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 74:21]
  assign io_out_valid = io_in_0_valid; // @[Arbiter.scala 55:16]
  assign io_out_bits_rd = io_in_0_bits_rd; // @[Arbiter.scala 56:15]
  assign io_out_bits_data = io_in_0_bits_data; // @[Arbiter.scala 56:15]
endmodule
module ComposerAcc(
  input          clock,
  input          reset,
  input          auto_EnergyCalc_memory_endpoint_identity_out_4_a_ready,
  output         auto_EnergyCalc_memory_endpoint_identity_out_4_a_valid,
  output [2:0]   auto_EnergyCalc_memory_endpoint_identity_out_4_a_bits_size,
  output [3:0]   auto_EnergyCalc_memory_endpoint_identity_out_4_a_bits_source,
  output [33:0]  auto_EnergyCalc_memory_endpoint_identity_out_4_a_bits_address,
  output [63:0]  auto_EnergyCalc_memory_endpoint_identity_out_4_a_bits_mask,
  output         auto_EnergyCalc_memory_endpoint_identity_out_4_d_ready,
  input          auto_EnergyCalc_memory_endpoint_identity_out_4_d_valid,
  input  [3:0]   auto_EnergyCalc_memory_endpoint_identity_out_4_d_bits_source,
  input          auto_EnergyCalc_memory_endpoint_identity_out_3_a_ready,
  output         auto_EnergyCalc_memory_endpoint_identity_out_3_a_valid,
  output [2:0]   auto_EnergyCalc_memory_endpoint_identity_out_3_a_bits_size,
  output [3:0]   auto_EnergyCalc_memory_endpoint_identity_out_3_a_bits_source,
  output [33:0]  auto_EnergyCalc_memory_endpoint_identity_out_3_a_bits_address,
  output [63:0]  auto_EnergyCalc_memory_endpoint_identity_out_3_a_bits_mask,
  output         auto_EnergyCalc_memory_endpoint_identity_out_3_d_ready,
  input          auto_EnergyCalc_memory_endpoint_identity_out_3_d_valid,
  input  [3:0]   auto_EnergyCalc_memory_endpoint_identity_out_3_d_bits_source,
  input          auto_EnergyCalc_memory_endpoint_identity_out_2_a_ready,
  output         auto_EnergyCalc_memory_endpoint_identity_out_2_a_valid,
  output [2:0]   auto_EnergyCalc_memory_endpoint_identity_out_2_a_bits_size,
  output [3:0]   auto_EnergyCalc_memory_endpoint_identity_out_2_a_bits_source,
  output [33:0]  auto_EnergyCalc_memory_endpoint_identity_out_2_a_bits_address,
  output [63:0]  auto_EnergyCalc_memory_endpoint_identity_out_2_a_bits_mask,
  output         auto_EnergyCalc_memory_endpoint_identity_out_2_d_ready,
  input          auto_EnergyCalc_memory_endpoint_identity_out_2_d_valid,
  input  [3:0]   auto_EnergyCalc_memory_endpoint_identity_out_2_d_bits_source,
  input          auto_EnergyCalc_memory_endpoint_identity_out_1_a_ready,
  output         auto_EnergyCalc_memory_endpoint_identity_out_1_a_valid,
  output [2:0]   auto_EnergyCalc_memory_endpoint_identity_out_1_a_bits_size,
  output [3:0]   auto_EnergyCalc_memory_endpoint_identity_out_1_a_bits_source,
  output [33:0]  auto_EnergyCalc_memory_endpoint_identity_out_1_a_bits_address,
  output [63:0]  auto_EnergyCalc_memory_endpoint_identity_out_1_a_bits_mask,
  output         auto_EnergyCalc_memory_endpoint_identity_out_1_d_ready,
  input          auto_EnergyCalc_memory_endpoint_identity_out_1_d_valid,
  input  [3:0]   auto_EnergyCalc_memory_endpoint_identity_out_1_d_bits_source,
  input  [511:0] auto_EnergyCalc_memory_endpoint_identity_out_1_d_bits_data,
  input          auto_EnergyCalc_memory_endpoint_identity_out_0_a_ready,
  output         auto_EnergyCalc_memory_endpoint_identity_out_0_a_valid,
  output         auto_EnergyCalc_memory_endpoint_identity_out_0_a_bits_source,
  output [33:0]  auto_EnergyCalc_memory_endpoint_identity_out_0_a_bits_address,
  output [63:0]  auto_EnergyCalc_memory_endpoint_identity_out_0_a_bits_mask,
  output [511:0] auto_EnergyCalc_memory_endpoint_identity_out_0_a_bits_data,
  output         auto_EnergyCalc_memory_endpoint_identity_out_0_d_ready,
  input          auto_EnergyCalc_memory_endpoint_identity_out_0_d_valid,
  input          auto_EnergyCalc_memory_endpoint_identity_out_0_d_bits_source,
  output         io_cmd_ready,
  input          io_cmd_valid,
  input  [6:0]   io_cmd_bits_inst_funct,
  input  [4:0]   io_cmd_bits_inst_rs2,
  input  [4:0]   io_cmd_bits_inst_rs1,
  input  [6:0]   io_cmd_bits_inst_opcode,
  input  [63:0]  io_cmd_bits_rs1,
  input  [63:0]  io_cmd_bits_rs2,
  input          io_resp_ready,
  output         io_resp_valid,
  output [4:0]   io_resp_bits_rd,
  output [63:0]  io_resp_bits_data
);
  wire  EnergyCalc_clock; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_reset; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_auto_memory_endpoint_identity_out_4_a_ready; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_auto_memory_endpoint_identity_out_4_a_valid; // @[Accelerator.scala 33:16]
  wire [2:0] EnergyCalc_auto_memory_endpoint_identity_out_4_a_bits_size; // @[Accelerator.scala 33:16]
  wire [3:0] EnergyCalc_auto_memory_endpoint_identity_out_4_a_bits_source; // @[Accelerator.scala 33:16]
  wire [33:0] EnergyCalc_auto_memory_endpoint_identity_out_4_a_bits_address; // @[Accelerator.scala 33:16]
  wire [63:0] EnergyCalc_auto_memory_endpoint_identity_out_4_a_bits_mask; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_auto_memory_endpoint_identity_out_4_d_ready; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_auto_memory_endpoint_identity_out_4_d_valid; // @[Accelerator.scala 33:16]
  wire [3:0] EnergyCalc_auto_memory_endpoint_identity_out_4_d_bits_source; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_auto_memory_endpoint_identity_out_3_a_ready; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_auto_memory_endpoint_identity_out_3_a_valid; // @[Accelerator.scala 33:16]
  wire [2:0] EnergyCalc_auto_memory_endpoint_identity_out_3_a_bits_size; // @[Accelerator.scala 33:16]
  wire [3:0] EnergyCalc_auto_memory_endpoint_identity_out_3_a_bits_source; // @[Accelerator.scala 33:16]
  wire [33:0] EnergyCalc_auto_memory_endpoint_identity_out_3_a_bits_address; // @[Accelerator.scala 33:16]
  wire [63:0] EnergyCalc_auto_memory_endpoint_identity_out_3_a_bits_mask; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_auto_memory_endpoint_identity_out_3_d_ready; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_auto_memory_endpoint_identity_out_3_d_valid; // @[Accelerator.scala 33:16]
  wire [3:0] EnergyCalc_auto_memory_endpoint_identity_out_3_d_bits_source; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_auto_memory_endpoint_identity_out_2_a_ready; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_auto_memory_endpoint_identity_out_2_a_valid; // @[Accelerator.scala 33:16]
  wire [2:0] EnergyCalc_auto_memory_endpoint_identity_out_2_a_bits_size; // @[Accelerator.scala 33:16]
  wire [3:0] EnergyCalc_auto_memory_endpoint_identity_out_2_a_bits_source; // @[Accelerator.scala 33:16]
  wire [33:0] EnergyCalc_auto_memory_endpoint_identity_out_2_a_bits_address; // @[Accelerator.scala 33:16]
  wire [63:0] EnergyCalc_auto_memory_endpoint_identity_out_2_a_bits_mask; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_auto_memory_endpoint_identity_out_2_d_ready; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_auto_memory_endpoint_identity_out_2_d_valid; // @[Accelerator.scala 33:16]
  wire [3:0] EnergyCalc_auto_memory_endpoint_identity_out_2_d_bits_source; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_auto_memory_endpoint_identity_out_1_a_ready; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_auto_memory_endpoint_identity_out_1_a_valid; // @[Accelerator.scala 33:16]
  wire [2:0] EnergyCalc_auto_memory_endpoint_identity_out_1_a_bits_size; // @[Accelerator.scala 33:16]
  wire [3:0] EnergyCalc_auto_memory_endpoint_identity_out_1_a_bits_source; // @[Accelerator.scala 33:16]
  wire [33:0] EnergyCalc_auto_memory_endpoint_identity_out_1_a_bits_address; // @[Accelerator.scala 33:16]
  wire [63:0] EnergyCalc_auto_memory_endpoint_identity_out_1_a_bits_mask; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_auto_memory_endpoint_identity_out_1_d_ready; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_auto_memory_endpoint_identity_out_1_d_valid; // @[Accelerator.scala 33:16]
  wire [3:0] EnergyCalc_auto_memory_endpoint_identity_out_1_d_bits_source; // @[Accelerator.scala 33:16]
  wire [511:0] EnergyCalc_auto_memory_endpoint_identity_out_1_d_bits_data; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_auto_memory_endpoint_identity_out_0_a_ready; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_auto_memory_endpoint_identity_out_0_a_valid; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_auto_memory_endpoint_identity_out_0_a_bits_source; // @[Accelerator.scala 33:16]
  wire [33:0] EnergyCalc_auto_memory_endpoint_identity_out_0_a_bits_address; // @[Accelerator.scala 33:16]
  wire [63:0] EnergyCalc_auto_memory_endpoint_identity_out_0_a_bits_mask; // @[Accelerator.scala 33:16]
  wire [511:0] EnergyCalc_auto_memory_endpoint_identity_out_0_a_bits_data; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_auto_memory_endpoint_identity_out_0_d_ready; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_auto_memory_endpoint_identity_out_0_d_valid; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_auto_memory_endpoint_identity_out_0_d_bits_source; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_sw_io_cmd_ready; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_sw_io_cmd_valid; // @[Accelerator.scala 33:16]
  wire [4:0] EnergyCalc_sw_io_cmd_bits_inst_rs1; // @[Accelerator.scala 33:16]
  wire [4:0] EnergyCalc_sw_io_cmd_bits_inst_rs2; // @[Accelerator.scala 33:16]
  wire [2:0] EnergyCalc_sw_io_cmd_bits_inst_funct; // @[Accelerator.scala 33:16]
  wire [7:0] EnergyCalc_sw_io_cmd_bits_core_id; // @[Accelerator.scala 33:16]
  wire [55:0] EnergyCalc_sw_io_cmd_bits_payload1; // @[Accelerator.scala 33:16]
  wire [63:0] EnergyCalc_sw_io_cmd_bits_payload2; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_sw_io_resp_ready; // @[Accelerator.scala 33:16]
  wire  EnergyCalc_sw_io_resp_valid; // @[Accelerator.scala 33:16]
  wire [4:0] EnergyCalc_sw_io_resp_bits_rd; // @[Accelerator.scala 33:16]
  wire [3:0] EnergyCalc_sw_io_resp_bits_system_id; // @[Accelerator.scala 33:16]
  wire [7:0] EnergyCalc_sw_io_resp_bits_core_id; // @[Accelerator.scala 33:16]
  wire [46:0] EnergyCalc_sw_io_resp_bits_data; // @[Accelerator.scala 33:16]
  wire  cmd_clock; // @[Decoupled.scala 375:21]
  wire  cmd_reset; // @[Decoupled.scala 375:21]
  wire  cmd_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  cmd_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [6:0] cmd_io_enq_bits_inst_funct; // @[Decoupled.scala 375:21]
  wire [4:0] cmd_io_enq_bits_inst_rs2; // @[Decoupled.scala 375:21]
  wire [4:0] cmd_io_enq_bits_inst_rs1; // @[Decoupled.scala 375:21]
  wire [6:0] cmd_io_enq_bits_inst_opcode; // @[Decoupled.scala 375:21]
  wire [63:0] cmd_io_enq_bits_rs1; // @[Decoupled.scala 375:21]
  wire [63:0] cmd_io_enq_bits_rs2; // @[Decoupled.scala 375:21]
  wire  cmd_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  cmd_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [6:0] cmd_io_deq_bits_inst_funct; // @[Decoupled.scala 375:21]
  wire [4:0] cmd_io_deq_bits_inst_rs2; // @[Decoupled.scala 375:21]
  wire [4:0] cmd_io_deq_bits_inst_rs1; // @[Decoupled.scala 375:21]
  wire [6:0] cmd_io_deq_bits_inst_opcode; // @[Decoupled.scala 375:21]
  wire [63:0] cmd_io_deq_bits_rs1; // @[Decoupled.scala 375:21]
  wire [63:0] cmd_io_deq_bits_rs2; // @[Decoupled.scala 375:21]
  wire  cmdArb_io_in_0_ready; // @[Accelerator.scala 63:22]
  wire  cmdArb_io_in_0_valid; // @[Accelerator.scala 63:22]
  wire [6:0] cmdArb_io_in_0_bits_inst_funct; // @[Accelerator.scala 63:22]
  wire [4:0] cmdArb_io_in_0_bits_inst_rs2; // @[Accelerator.scala 63:22]
  wire [4:0] cmdArb_io_in_0_bits_inst_rs1; // @[Accelerator.scala 63:22]
  wire [6:0] cmdArb_io_in_0_bits_inst_opcode; // @[Accelerator.scala 63:22]
  wire [63:0] cmdArb_io_in_0_bits_rs1; // @[Accelerator.scala 63:22]
  wire [63:0] cmdArb_io_in_0_bits_rs2; // @[Accelerator.scala 63:22]
  wire  cmdArb_io_out_ready; // @[Accelerator.scala 63:22]
  wire  cmdArb_io_out_valid; // @[Accelerator.scala 63:22]
  wire [6:0] cmdArb_io_out_bits_inst_funct; // @[Accelerator.scala 63:22]
  wire [4:0] cmdArb_io_out_bits_inst_rs2; // @[Accelerator.scala 63:22]
  wire [4:0] cmdArb_io_out_bits_inst_rs1; // @[Accelerator.scala 63:22]
  wire [6:0] cmdArb_io_out_bits_inst_opcode; // @[Accelerator.scala 63:22]
  wire [63:0] cmdArb_io_out_bits_rs1; // @[Accelerator.scala 63:22]
  wire [63:0] cmdArb_io_out_bits_rs2; // @[Accelerator.scala 63:22]
  wire  cmdRouter_clock; // @[Accelerator.scala 69:25]
  wire  cmdRouter_reset; // @[Accelerator.scala 69:25]
  wire  cmdRouter_io_in_ready; // @[Accelerator.scala 69:25]
  wire  cmdRouter_io_in_valid; // @[Accelerator.scala 69:25]
  wire [6:0] cmdRouter_io_in_bits_inst_funct; // @[Accelerator.scala 69:25]
  wire [4:0] cmdRouter_io_in_bits_inst_rs2; // @[Accelerator.scala 69:25]
  wire [4:0] cmdRouter_io_in_bits_inst_rs1; // @[Accelerator.scala 69:25]
  wire [6:0] cmdRouter_io_in_bits_inst_opcode; // @[Accelerator.scala 69:25]
  wire [63:0] cmdRouter_io_in_bits_rs1; // @[Accelerator.scala 69:25]
  wire [63:0] cmdRouter_io_in_bits_rs2; // @[Accelerator.scala 69:25]
  wire  cmdRouter_io_out_0_ready; // @[Accelerator.scala 69:25]
  wire  cmdRouter_io_out_0_valid; // @[Accelerator.scala 69:25]
  wire  cmdRouter_io_out_1_ready; // @[Accelerator.scala 69:25]
  wire  cmdRouter_io_out_1_valid; // @[Accelerator.scala 69:25]
  wire [6:0] cmdRouter_io_out_1_bits_inst_funct; // @[Accelerator.scala 69:25]
  wire [4:0] cmdRouter_io_out_1_bits_inst_rs2; // @[Accelerator.scala 69:25]
  wire [4:0] cmdRouter_io_out_1_bits_inst_rs1; // @[Accelerator.scala 69:25]
  wire [63:0] cmdRouter_io_out_1_bits_rs1; // @[Accelerator.scala 69:25]
  wire [63:0] cmdRouter_io_out_1_bits_rs2; // @[Accelerator.scala 69:25]
  wire
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_clock
    ; // @[Accelerator.scala 100:27]
  wire
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_reset
    ; // @[Accelerator.scala 100:27]
  wire
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_enq_ready
    ; // @[Accelerator.scala 100:27]
  wire
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_enq_valid
    ; // @[Accelerator.scala 100:27]
  wire [4:0]
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_enq_bits_inst_rs1
    ; // @[Accelerator.scala 100:27]
  wire [4:0]
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_enq_bits_inst_rs2
    ; // @[Accelerator.scala 100:27]
  wire [2:0]
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_enq_bits_inst_funct
    ; // @[Accelerator.scala 100:27]
  wire [7:0]
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_enq_bits_core_id
    ; // @[Accelerator.scala 100:27]
  wire [55:0]
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_enq_bits_payload1
    ; // @[Accelerator.scala 100:27]
  wire [63:0]
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_enq_bits_payload2
    ; // @[Accelerator.scala 100:27]
  wire
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_deq_ready
    ; // @[Accelerator.scala 100:27]
  wire
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_deq_valid
    ; // @[Accelerator.scala 100:27]
  wire [4:0]
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_deq_bits_inst_rs1
    ; // @[Accelerator.scala 100:27]
  wire [4:0]
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_deq_bits_inst_rs2
    ; // @[Accelerator.scala 100:27]
  wire [2:0]
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_deq_bits_inst_funct
    ; // @[Accelerator.scala 100:27]
  wire [7:0]
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_deq_bits_core_id
    ; // @[Accelerator.scala 100:27]
  wire [55:0]
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_deq_bits_payload1
    ; // @[Accelerator.scala 100:27]
  wire [63:0]
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_deq_bits_payload2
    ; // @[Accelerator.scala 100:27]
  wire  respArbiter_io_in_0_ready; // @[Accelerator.scala 127:29]
  wire  respArbiter_io_in_0_valid; // @[Accelerator.scala 127:29]
  wire [4:0] respArbiter_io_in_0_bits_rd; // @[Accelerator.scala 127:29]
  wire [63:0] respArbiter_io_in_0_bits_data; // @[Accelerator.scala 127:29]
  wire  respArbiter_io_out_ready; // @[Accelerator.scala 127:29]
  wire  respArbiter_io_out_valid; // @[Accelerator.scala 127:29]
  wire [4:0] respArbiter_io_out_bits_rd; // @[Accelerator.scala 127:29]
  wire [63:0] respArbiter_io_out_bits_data; // @[Accelerator.scala 127:29]
  wire [3:0] accCmd_bits_inst_system_id = cmdRouter_io_out_1_bits_inst_funct[6:3]; // @[Accelerator.scala 84:68]
  reg  waitingToFlush; // @[Accelerator.scala 93:31]
  wire  _T = cmdRouter_io_out_0_ready & cmdRouter_io_out_0_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_0 = _T | waitingToFlush; // @[Accelerator.scala 95:35 96:20 93:31]
  wire  accCmd_valid = cmdRouter_io_out_1_valid; // @[Accelerator.scala 72:20 73:16]
  wire [51:0] respArbiter_io_in_0_bits_data_lo = {EnergyCalc_sw_io_resp_bits_rd,EnergyCalc_sw_io_resp_bits_data}; // @[Cat.scala 33:92]
  wire [11:0] respArbiter_io_in_0_bits_data_hi = {EnergyCalc_sw_io_resp_bits_system_id,
    EnergyCalc_sw_io_resp_bits_core_id}; // @[Cat.scala 33:92]
  ComposerSystem EnergyCalc ( // @[Accelerator.scala 33:16]
    .clock(EnergyCalc_clock),
    .reset(EnergyCalc_reset),
    .auto_memory_endpoint_identity_out_4_a_ready(EnergyCalc_auto_memory_endpoint_identity_out_4_a_ready),
    .auto_memory_endpoint_identity_out_4_a_valid(EnergyCalc_auto_memory_endpoint_identity_out_4_a_valid),
    .auto_memory_endpoint_identity_out_4_a_bits_size(EnergyCalc_auto_memory_endpoint_identity_out_4_a_bits_size),
    .auto_memory_endpoint_identity_out_4_a_bits_source(EnergyCalc_auto_memory_endpoint_identity_out_4_a_bits_source),
    .auto_memory_endpoint_identity_out_4_a_bits_address(EnergyCalc_auto_memory_endpoint_identity_out_4_a_bits_address),
    .auto_memory_endpoint_identity_out_4_a_bits_mask(EnergyCalc_auto_memory_endpoint_identity_out_4_a_bits_mask),
    .auto_memory_endpoint_identity_out_4_d_ready(EnergyCalc_auto_memory_endpoint_identity_out_4_d_ready),
    .auto_memory_endpoint_identity_out_4_d_valid(EnergyCalc_auto_memory_endpoint_identity_out_4_d_valid),
    .auto_memory_endpoint_identity_out_4_d_bits_source(EnergyCalc_auto_memory_endpoint_identity_out_4_d_bits_source),
    .auto_memory_endpoint_identity_out_3_a_ready(EnergyCalc_auto_memory_endpoint_identity_out_3_a_ready),
    .auto_memory_endpoint_identity_out_3_a_valid(EnergyCalc_auto_memory_endpoint_identity_out_3_a_valid),
    .auto_memory_endpoint_identity_out_3_a_bits_size(EnergyCalc_auto_memory_endpoint_identity_out_3_a_bits_size),
    .auto_memory_endpoint_identity_out_3_a_bits_source(EnergyCalc_auto_memory_endpoint_identity_out_3_a_bits_source),
    .auto_memory_endpoint_identity_out_3_a_bits_address(EnergyCalc_auto_memory_endpoint_identity_out_3_a_bits_address),
    .auto_memory_endpoint_identity_out_3_a_bits_mask(EnergyCalc_auto_memory_endpoint_identity_out_3_a_bits_mask),
    .auto_memory_endpoint_identity_out_3_d_ready(EnergyCalc_auto_memory_endpoint_identity_out_3_d_ready),
    .auto_memory_endpoint_identity_out_3_d_valid(EnergyCalc_auto_memory_endpoint_identity_out_3_d_valid),
    .auto_memory_endpoint_identity_out_3_d_bits_source(EnergyCalc_auto_memory_endpoint_identity_out_3_d_bits_source),
    .auto_memory_endpoint_identity_out_2_a_ready(EnergyCalc_auto_memory_endpoint_identity_out_2_a_ready),
    .auto_memory_endpoint_identity_out_2_a_valid(EnergyCalc_auto_memory_endpoint_identity_out_2_a_valid),
    .auto_memory_endpoint_identity_out_2_a_bits_size(EnergyCalc_auto_memory_endpoint_identity_out_2_a_bits_size),
    .auto_memory_endpoint_identity_out_2_a_bits_source(EnergyCalc_auto_memory_endpoint_identity_out_2_a_bits_source),
    .auto_memory_endpoint_identity_out_2_a_bits_address(EnergyCalc_auto_memory_endpoint_identity_out_2_a_bits_address),
    .auto_memory_endpoint_identity_out_2_a_bits_mask(EnergyCalc_auto_memory_endpoint_identity_out_2_a_bits_mask),
    .auto_memory_endpoint_identity_out_2_d_ready(EnergyCalc_auto_memory_endpoint_identity_out_2_d_ready),
    .auto_memory_endpoint_identity_out_2_d_valid(EnergyCalc_auto_memory_endpoint_identity_out_2_d_valid),
    .auto_memory_endpoint_identity_out_2_d_bits_source(EnergyCalc_auto_memory_endpoint_identity_out_2_d_bits_source),
    .auto_memory_endpoint_identity_out_1_a_ready(EnergyCalc_auto_memory_endpoint_identity_out_1_a_ready),
    .auto_memory_endpoint_identity_out_1_a_valid(EnergyCalc_auto_memory_endpoint_identity_out_1_a_valid),
    .auto_memory_endpoint_identity_out_1_a_bits_size(EnergyCalc_auto_memory_endpoint_identity_out_1_a_bits_size),
    .auto_memory_endpoint_identity_out_1_a_bits_source(EnergyCalc_auto_memory_endpoint_identity_out_1_a_bits_source),
    .auto_memory_endpoint_identity_out_1_a_bits_address(EnergyCalc_auto_memory_endpoint_identity_out_1_a_bits_address),
    .auto_memory_endpoint_identity_out_1_a_bits_mask(EnergyCalc_auto_memory_endpoint_identity_out_1_a_bits_mask),
    .auto_memory_endpoint_identity_out_1_d_ready(EnergyCalc_auto_memory_endpoint_identity_out_1_d_ready),
    .auto_memory_endpoint_identity_out_1_d_valid(EnergyCalc_auto_memory_endpoint_identity_out_1_d_valid),
    .auto_memory_endpoint_identity_out_1_d_bits_source(EnergyCalc_auto_memory_endpoint_identity_out_1_d_bits_source),
    .auto_memory_endpoint_identity_out_1_d_bits_data(EnergyCalc_auto_memory_endpoint_identity_out_1_d_bits_data),
    .auto_memory_endpoint_identity_out_0_a_ready(EnergyCalc_auto_memory_endpoint_identity_out_0_a_ready),
    .auto_memory_endpoint_identity_out_0_a_valid(EnergyCalc_auto_memory_endpoint_identity_out_0_a_valid),
    .auto_memory_endpoint_identity_out_0_a_bits_source(EnergyCalc_auto_memory_endpoint_identity_out_0_a_bits_source),
    .auto_memory_endpoint_identity_out_0_a_bits_address(EnergyCalc_auto_memory_endpoint_identity_out_0_a_bits_address),
    .auto_memory_endpoint_identity_out_0_a_bits_mask(EnergyCalc_auto_memory_endpoint_identity_out_0_a_bits_mask),
    .auto_memory_endpoint_identity_out_0_a_bits_data(EnergyCalc_auto_memory_endpoint_identity_out_0_a_bits_data),
    .auto_memory_endpoint_identity_out_0_d_ready(EnergyCalc_auto_memory_endpoint_identity_out_0_d_ready),
    .auto_memory_endpoint_identity_out_0_d_valid(EnergyCalc_auto_memory_endpoint_identity_out_0_d_valid),
    .auto_memory_endpoint_identity_out_0_d_bits_source(EnergyCalc_auto_memory_endpoint_identity_out_0_d_bits_source),
    .sw_io_cmd_ready(EnergyCalc_sw_io_cmd_ready),
    .sw_io_cmd_valid(EnergyCalc_sw_io_cmd_valid),
    .sw_io_cmd_bits_inst_rs1(EnergyCalc_sw_io_cmd_bits_inst_rs1),
    .sw_io_cmd_bits_inst_rs2(EnergyCalc_sw_io_cmd_bits_inst_rs2),
    .sw_io_cmd_bits_inst_funct(EnergyCalc_sw_io_cmd_bits_inst_funct),
    .sw_io_cmd_bits_core_id(EnergyCalc_sw_io_cmd_bits_core_id),
    .sw_io_cmd_bits_payload1(EnergyCalc_sw_io_cmd_bits_payload1),
    .sw_io_cmd_bits_payload2(EnergyCalc_sw_io_cmd_bits_payload2),
    .sw_io_resp_ready(EnergyCalc_sw_io_resp_ready),
    .sw_io_resp_valid(EnergyCalc_sw_io_resp_valid),
    .sw_io_resp_bits_rd(EnergyCalc_sw_io_resp_bits_rd),
    .sw_io_resp_bits_system_id(EnergyCalc_sw_io_resp_bits_system_id),
    .sw_io_resp_bits_core_id(EnergyCalc_sw_io_resp_bits_core_id),
    .sw_io_resp_bits_data(EnergyCalc_sw_io_resp_bits_data)
  );
  Queue_3 cmd ( // @[Decoupled.scala 375:21]
    .clock(cmd_clock),
    .reset(cmd_reset),
    .io_enq_ready(cmd_io_enq_ready),
    .io_enq_valid(cmd_io_enq_valid),
    .io_enq_bits_inst_funct(cmd_io_enq_bits_inst_funct),
    .io_enq_bits_inst_rs2(cmd_io_enq_bits_inst_rs2),
    .io_enq_bits_inst_rs1(cmd_io_enq_bits_inst_rs1),
    .io_enq_bits_inst_opcode(cmd_io_enq_bits_inst_opcode),
    .io_enq_bits_rs1(cmd_io_enq_bits_rs1),
    .io_enq_bits_rs2(cmd_io_enq_bits_rs2),
    .io_deq_ready(cmd_io_deq_ready),
    .io_deq_valid(cmd_io_deq_valid),
    .io_deq_bits_inst_funct(cmd_io_deq_bits_inst_funct),
    .io_deq_bits_inst_rs2(cmd_io_deq_bits_inst_rs2),
    .io_deq_bits_inst_rs1(cmd_io_deq_bits_inst_rs1),
    .io_deq_bits_inst_opcode(cmd_io_deq_bits_inst_opcode),
    .io_deq_bits_rs1(cmd_io_deq_bits_rs1),
    .io_deq_bits_rs2(cmd_io_deq_bits_rs2)
  );
  RRArbiter_1 cmdArb ( // @[Accelerator.scala 63:22]
    .io_in_0_ready(cmdArb_io_in_0_ready),
    .io_in_0_valid(cmdArb_io_in_0_valid),
    .io_in_0_bits_inst_funct(cmdArb_io_in_0_bits_inst_funct),
    .io_in_0_bits_inst_rs2(cmdArb_io_in_0_bits_inst_rs2),
    .io_in_0_bits_inst_rs1(cmdArb_io_in_0_bits_inst_rs1),
    .io_in_0_bits_inst_opcode(cmdArb_io_in_0_bits_inst_opcode),
    .io_in_0_bits_rs1(cmdArb_io_in_0_bits_rs1),
    .io_in_0_bits_rs2(cmdArb_io_in_0_bits_rs2),
    .io_out_ready(cmdArb_io_out_ready),
    .io_out_valid(cmdArb_io_out_valid),
    .io_out_bits_inst_funct(cmdArb_io_out_bits_inst_funct),
    .io_out_bits_inst_rs2(cmdArb_io_out_bits_inst_rs2),
    .io_out_bits_inst_rs1(cmdArb_io_out_bits_inst_rs1),
    .io_out_bits_inst_opcode(cmdArb_io_out_bits_inst_opcode),
    .io_out_bits_rs1(cmdArb_io_out_bits_rs1),
    .io_out_bits_rs2(cmdArb_io_out_bits_rs2)
  );
  RoccCommandRouter cmdRouter ( // @[Accelerator.scala 69:25]
    .clock(cmdRouter_clock),
    .reset(cmdRouter_reset),
    .io_in_ready(cmdRouter_io_in_ready),
    .io_in_valid(cmdRouter_io_in_valid),
    .io_in_bits_inst_funct(cmdRouter_io_in_bits_inst_funct),
    .io_in_bits_inst_rs2(cmdRouter_io_in_bits_inst_rs2),
    .io_in_bits_inst_rs1(cmdRouter_io_in_bits_inst_rs1),
    .io_in_bits_inst_opcode(cmdRouter_io_in_bits_inst_opcode),
    .io_in_bits_rs1(cmdRouter_io_in_bits_rs1),
    .io_in_bits_rs2(cmdRouter_io_in_bits_rs2),
    .io_out_0_ready(cmdRouter_io_out_0_ready),
    .io_out_0_valid(cmdRouter_io_out_0_valid),
    .io_out_1_ready(cmdRouter_io_out_1_ready),
    .io_out_1_valid(cmdRouter_io_out_1_valid),
    .io_out_1_bits_inst_funct(cmdRouter_io_out_1_bits_inst_funct),
    .io_out_1_bits_inst_rs2(cmdRouter_io_out_1_bits_inst_rs2),
    .io_out_1_bits_inst_rs1(cmdRouter_io_out_1_bits_inst_rs1),
    .io_out_1_bits_rs1(cmdRouter_io_out_1_bits_rs1),
    .io_out_1_bits_rs2(cmdRouter_io_out_1_bits_rs2)
  );
  Queue
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue
     ( // @[Accelerator.scala 100:27]
    .clock(
      systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_clock
      ),
    .reset(
      systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_reset
      ),
    .io_enq_ready(
      systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_enq_ready
      ),
    .io_enq_valid(
      systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_enq_valid
      ),
    .io_enq_bits_inst_rs1(
      systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_enq_bits_inst_rs1
      ),
    .io_enq_bits_inst_rs2(
      systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_enq_bits_inst_rs2
      ),
    .io_enq_bits_inst_funct(
      systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_enq_bits_inst_funct
      ),
    .io_enq_bits_core_id(
      systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_enq_bits_core_id
      ),
    .io_enq_bits_payload1(
      systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_enq_bits_payload1
      ),
    .io_enq_bits_payload2(
      systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_enq_bits_payload2
      ),
    .io_deq_ready(
      systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_deq_ready
      ),
    .io_deq_valid(
      systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_deq_valid
      ),
    .io_deq_bits_inst_rs1(
      systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_deq_bits_inst_rs1
      ),
    .io_deq_bits_inst_rs2(
      systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_deq_bits_inst_rs2
      ),
    .io_deq_bits_inst_funct(
      systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_deq_bits_inst_funct
      ),
    .io_deq_bits_core_id(
      systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_deq_bits_core_id
      ),
    .io_deq_bits_payload1(
      systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_deq_bits_payload1
      ),
    .io_deq_bits_payload2(
      systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_deq_bits_payload2
      )
  );
  RRArbiter_2 respArbiter ( // @[Accelerator.scala 127:29]
    .io_in_0_ready(respArbiter_io_in_0_ready),
    .io_in_0_valid(respArbiter_io_in_0_valid),
    .io_in_0_bits_rd(respArbiter_io_in_0_bits_rd),
    .io_in_0_bits_data(respArbiter_io_in_0_bits_data),
    .io_out_ready(respArbiter_io_out_ready),
    .io_out_valid(respArbiter_io_out_valid),
    .io_out_bits_rd(respArbiter_io_out_bits_rd),
    .io_out_bits_data(respArbiter_io_out_bits_data)
  );
  assign auto_EnergyCalc_memory_endpoint_identity_out_4_a_valid = EnergyCalc_auto_memory_endpoint_identity_out_4_a_valid
    ; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_4_a_bits_size =
    EnergyCalc_auto_memory_endpoint_identity_out_4_a_bits_size; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_4_a_bits_source =
    EnergyCalc_auto_memory_endpoint_identity_out_4_a_bits_source; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_4_a_bits_address =
    EnergyCalc_auto_memory_endpoint_identity_out_4_a_bits_address; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_4_a_bits_mask =
    EnergyCalc_auto_memory_endpoint_identity_out_4_a_bits_mask; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_4_d_ready = EnergyCalc_auto_memory_endpoint_identity_out_4_d_ready
    ; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_3_a_valid = EnergyCalc_auto_memory_endpoint_identity_out_3_a_valid
    ; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_3_a_bits_size =
    EnergyCalc_auto_memory_endpoint_identity_out_3_a_bits_size; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_3_a_bits_source =
    EnergyCalc_auto_memory_endpoint_identity_out_3_a_bits_source; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_3_a_bits_address =
    EnergyCalc_auto_memory_endpoint_identity_out_3_a_bits_address; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_3_a_bits_mask =
    EnergyCalc_auto_memory_endpoint_identity_out_3_a_bits_mask; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_3_d_ready = EnergyCalc_auto_memory_endpoint_identity_out_3_d_ready
    ; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_2_a_valid = EnergyCalc_auto_memory_endpoint_identity_out_2_a_valid
    ; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_2_a_bits_size =
    EnergyCalc_auto_memory_endpoint_identity_out_2_a_bits_size; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_2_a_bits_source =
    EnergyCalc_auto_memory_endpoint_identity_out_2_a_bits_source; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_2_a_bits_address =
    EnergyCalc_auto_memory_endpoint_identity_out_2_a_bits_address; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_2_a_bits_mask =
    EnergyCalc_auto_memory_endpoint_identity_out_2_a_bits_mask; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_2_d_ready = EnergyCalc_auto_memory_endpoint_identity_out_2_d_ready
    ; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_1_a_valid = EnergyCalc_auto_memory_endpoint_identity_out_1_a_valid
    ; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_1_a_bits_size =
    EnergyCalc_auto_memory_endpoint_identity_out_1_a_bits_size; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_1_a_bits_source =
    EnergyCalc_auto_memory_endpoint_identity_out_1_a_bits_source; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_1_a_bits_address =
    EnergyCalc_auto_memory_endpoint_identity_out_1_a_bits_address; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_1_a_bits_mask =
    EnergyCalc_auto_memory_endpoint_identity_out_1_a_bits_mask; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_1_d_ready = EnergyCalc_auto_memory_endpoint_identity_out_1_d_ready
    ; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_0_a_valid = EnergyCalc_auto_memory_endpoint_identity_out_0_a_valid
    ; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_0_a_bits_source =
    EnergyCalc_auto_memory_endpoint_identity_out_0_a_bits_source; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_0_a_bits_address =
    EnergyCalc_auto_memory_endpoint_identity_out_0_a_bits_address; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_0_a_bits_mask =
    EnergyCalc_auto_memory_endpoint_identity_out_0_a_bits_mask; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_0_a_bits_data =
    EnergyCalc_auto_memory_endpoint_identity_out_0_a_bits_data; // @[LazyModule.scala 368:12]
  assign auto_EnergyCalc_memory_endpoint_identity_out_0_d_ready = EnergyCalc_auto_memory_endpoint_identity_out_0_d_ready
    ; // @[LazyModule.scala 368:12]
  assign io_cmd_ready = cmd_io_enq_ready; // @[Decoupled.scala 379:17]
  assign io_resp_valid = respArbiter_io_out_valid; // @[Accelerator.scala 134:24]
  assign io_resp_bits_rd = respArbiter_io_out_bits_rd; // @[Accelerator.scala 134:24]
  assign io_resp_bits_data = respArbiter_io_out_bits_data; // @[Accelerator.scala 134:24]
  assign EnergyCalc_clock = clock;
  assign EnergyCalc_reset = reset;
  assign EnergyCalc_auto_memory_endpoint_identity_out_4_a_ready = auto_EnergyCalc_memory_endpoint_identity_out_4_a_ready
    ; // @[LazyModule.scala 368:12]
  assign EnergyCalc_auto_memory_endpoint_identity_out_4_d_valid = auto_EnergyCalc_memory_endpoint_identity_out_4_d_valid
    ; // @[LazyModule.scala 368:12]
  assign EnergyCalc_auto_memory_endpoint_identity_out_4_d_bits_source =
    auto_EnergyCalc_memory_endpoint_identity_out_4_d_bits_source; // @[LazyModule.scala 368:12]
  assign EnergyCalc_auto_memory_endpoint_identity_out_3_a_ready = auto_EnergyCalc_memory_endpoint_identity_out_3_a_ready
    ; // @[LazyModule.scala 368:12]
  assign EnergyCalc_auto_memory_endpoint_identity_out_3_d_valid = auto_EnergyCalc_memory_endpoint_identity_out_3_d_valid
    ; // @[LazyModule.scala 368:12]
  assign EnergyCalc_auto_memory_endpoint_identity_out_3_d_bits_source =
    auto_EnergyCalc_memory_endpoint_identity_out_3_d_bits_source; // @[LazyModule.scala 368:12]
  assign EnergyCalc_auto_memory_endpoint_identity_out_2_a_ready = auto_EnergyCalc_memory_endpoint_identity_out_2_a_ready
    ; // @[LazyModule.scala 368:12]
  assign EnergyCalc_auto_memory_endpoint_identity_out_2_d_valid = auto_EnergyCalc_memory_endpoint_identity_out_2_d_valid
    ; // @[LazyModule.scala 368:12]
  assign EnergyCalc_auto_memory_endpoint_identity_out_2_d_bits_source =
    auto_EnergyCalc_memory_endpoint_identity_out_2_d_bits_source; // @[LazyModule.scala 368:12]
  assign EnergyCalc_auto_memory_endpoint_identity_out_1_a_ready = auto_EnergyCalc_memory_endpoint_identity_out_1_a_ready
    ; // @[LazyModule.scala 368:12]
  assign EnergyCalc_auto_memory_endpoint_identity_out_1_d_valid = auto_EnergyCalc_memory_endpoint_identity_out_1_d_valid
    ; // @[LazyModule.scala 368:12]
  assign EnergyCalc_auto_memory_endpoint_identity_out_1_d_bits_source =
    auto_EnergyCalc_memory_endpoint_identity_out_1_d_bits_source; // @[LazyModule.scala 368:12]
  assign EnergyCalc_auto_memory_endpoint_identity_out_1_d_bits_data =
    auto_EnergyCalc_memory_endpoint_identity_out_1_d_bits_data; // @[LazyModule.scala 368:12]
  assign EnergyCalc_auto_memory_endpoint_identity_out_0_a_ready = auto_EnergyCalc_memory_endpoint_identity_out_0_a_ready
    ; // @[LazyModule.scala 368:12]
  assign EnergyCalc_auto_memory_endpoint_identity_out_0_d_valid = auto_EnergyCalc_memory_endpoint_identity_out_0_d_valid
    ; // @[LazyModule.scala 368:12]
  assign EnergyCalc_auto_memory_endpoint_identity_out_0_d_bits_source =
    auto_EnergyCalc_memory_endpoint_identity_out_0_d_bits_source; // @[LazyModule.scala 368:12]
  assign EnergyCalc_sw_io_cmd_valid = waitingToFlush ? 1'h0 :
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_deq_valid
    ; // @[Accelerator.scala 116:26 113:37 118:45]
  assign EnergyCalc_sw_io_cmd_bits_inst_rs1 =
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_deq_bits_inst_rs1
    ; // @[Accelerator.scala 113:37]
  assign EnergyCalc_sw_io_cmd_bits_inst_rs2 =
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_deq_bits_inst_rs2
    ; // @[Accelerator.scala 113:37]
  assign EnergyCalc_sw_io_cmd_bits_inst_funct =
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_deq_bits_inst_funct
    ; // @[Accelerator.scala 113:37]
  assign EnergyCalc_sw_io_cmd_bits_core_id =
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_deq_bits_core_id
    ; // @[Accelerator.scala 113:37]
  assign EnergyCalc_sw_io_cmd_bits_payload1 =
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_deq_bits_payload1
    ; // @[Accelerator.scala 113:37]
  assign EnergyCalc_sw_io_cmd_bits_payload2 =
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_deq_bits_payload2
    ; // @[Accelerator.scala 113:37]
  assign EnergyCalc_sw_io_resp_ready = respArbiter_io_in_0_ready; // @[Accelerator.scala 132:19]
  assign cmd_clock = clock;
  assign cmd_reset = reset;
  assign cmd_io_enq_valid = io_cmd_valid; // @[Decoupled.scala 377:22]
  assign cmd_io_enq_bits_inst_funct = io_cmd_bits_inst_funct; // @[Decoupled.scala 378:21]
  assign cmd_io_enq_bits_inst_rs2 = io_cmd_bits_inst_rs2; // @[Decoupled.scala 378:21]
  assign cmd_io_enq_bits_inst_rs1 = io_cmd_bits_inst_rs1; // @[Decoupled.scala 378:21]
  assign cmd_io_enq_bits_inst_opcode = io_cmd_bits_inst_opcode; // @[Decoupled.scala 378:21]
  assign cmd_io_enq_bits_rs1 = io_cmd_bits_rs1; // @[Decoupled.scala 378:21]
  assign cmd_io_enq_bits_rs2 = io_cmd_bits_rs2; // @[Decoupled.scala 378:21]
  assign cmd_io_deq_ready = cmdArb_io_in_0_ready; // @[Accelerator.scala 64:19]
  assign cmdArb_io_in_0_valid = cmd_io_deq_valid; // @[Accelerator.scala 64:19]
  assign cmdArb_io_in_0_bits_inst_funct = cmd_io_deq_bits_inst_funct; // @[Accelerator.scala 64:19]
  assign cmdArb_io_in_0_bits_inst_rs2 = cmd_io_deq_bits_inst_rs2; // @[Accelerator.scala 64:19]
  assign cmdArb_io_in_0_bits_inst_rs1 = cmd_io_deq_bits_inst_rs1; // @[Accelerator.scala 64:19]
  assign cmdArb_io_in_0_bits_inst_opcode = cmd_io_deq_bits_inst_opcode; // @[Accelerator.scala 64:19]
  assign cmdArb_io_in_0_bits_rs1 = cmd_io_deq_bits_rs1; // @[Accelerator.scala 64:19]
  assign cmdArb_io_in_0_bits_rs2 = cmd_io_deq_bits_rs2; // @[Accelerator.scala 64:19]
  assign cmdArb_io_out_ready = cmdRouter_io_in_ready; // @[Accelerator.scala 70:19]
  assign cmdRouter_clock = clock;
  assign cmdRouter_reset = reset;
  assign cmdRouter_io_in_valid = cmdArb_io_out_valid; // @[Accelerator.scala 70:19]
  assign cmdRouter_io_in_bits_inst_funct = cmdArb_io_out_bits_inst_funct; // @[Accelerator.scala 70:19]
  assign cmdRouter_io_in_bits_inst_rs2 = cmdArb_io_out_bits_inst_rs2; // @[Accelerator.scala 70:19]
  assign cmdRouter_io_in_bits_inst_rs1 = cmdArb_io_out_bits_inst_rs1; // @[Accelerator.scala 70:19]
  assign cmdRouter_io_in_bits_inst_opcode = cmdArb_io_out_bits_inst_opcode; // @[Accelerator.scala 70:19]
  assign cmdRouter_io_in_bits_rs1 = cmdArb_io_out_bits_rs1; // @[Accelerator.scala 70:19]
  assign cmdRouter_io_in_bits_rs2 = cmdArb_io_out_bits_rs2; // @[Accelerator.scala 70:19]
  assign cmdRouter_io_out_0_ready = ~waitingToFlush; // @[Accelerator.scala 94:32]
  assign cmdRouter_io_out_1_ready = accCmd_bits_inst_system_id == 4'h0 &
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_enq_ready
    ; // @[Accelerator.scala 108:36 109:20 91:16]
  assign
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_clock
     = clock;
  assign
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_reset
     = reset;
  assign
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_enq_valid
     = accCmd_valid & 4'h0 == accCmd_bits_inst_system_id; // @[Accelerator.scala 106:44]
  assign
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_enq_bits_inst_rs1
     = cmdRouter_io_out_1_bits_inst_rs1; // @[Accelerator.scala 72:20 75:24]
  assign
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_enq_bits_inst_rs2
     = cmdRouter_io_out_1_bits_inst_rs2; // @[Accelerator.scala 72:20 76:24]
  assign
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_enq_bits_inst_funct
     = cmdRouter_io_out_1_bits_inst_funct[2:0]; // @[Accelerator.scala 83:64]
  assign
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_enq_bits_core_id
     = cmdRouter_io_out_1_bits_rs1[63:56]; // @[Accelerator.scala 86:54]
  assign
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_enq_bits_payload1
     = cmdRouter_io_out_1_bits_rs1[55:0]; // @[Accelerator.scala 87:55]
  assign
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_enq_bits_payload2
     = cmdRouter_io_out_1_bits_rs2; // @[Accelerator.scala 72:20 88:24]
  assign
    systemSoftwareResps_ComposerSystemParams1EnergyCalcdesignenergyCalcwithEnergyCalcanonfunlessinitgreater1anonfunapply1Lambda60810x0000000802076e905299be2bComposerCoreParamsListCChannelParamsWriteChannel1WriteChannelCChannelParamsdata1ScratchpadCChannelParamshalfNonBonded1ScratchpadCChannelParamsnonBonded1ScratchpadCChannelParamssolvated1Scratchpad00132truefalse_command_queue_io_deq_ready
     = waitingToFlush ? 1'h0 : EnergyCalc_sw_io_cmd_ready; // @[Accelerator.scala 116:26 117:30 113:37]
  assign respArbiter_io_in_0_valid = EnergyCalc_sw_io_resp_valid; // @[Accelerator.scala 131:19]
  assign respArbiter_io_in_0_bits_rd = EnergyCalc_sw_io_resp_bits_rd; // @[Accelerator.scala 130:21]
  assign respArbiter_io_in_0_bits_data = {respArbiter_io_in_0_bits_data_hi,respArbiter_io_in_0_bits_data_lo}; // @[Cat.scala 33:92]
  assign respArbiter_io_out_ready = io_resp_ready; // @[Accelerator.scala 134:24]
  always @(posedge clock) begin
    if (reset) begin // @[Accelerator.scala 93:31]
      waitingToFlush <= 1'h0; // @[Accelerator.scala 93:31]
    end else begin
      waitingToFlush <= _GEN_0;
    end
  end
endmodule
module TLXbar(
  input          clock,
  input          reset,
  output         auto_in_4_a_ready,
  input          auto_in_4_a_valid,
  input  [2:0]   auto_in_4_a_bits_size,
  input  [3:0]   auto_in_4_a_bits_source,
  input  [33:0]  auto_in_4_a_bits_address,
  input  [63:0]  auto_in_4_a_bits_mask,
  input          auto_in_4_d_ready,
  output         auto_in_4_d_valid,
  output [3:0]   auto_in_4_d_bits_source,
  output         auto_in_3_a_ready,
  input          auto_in_3_a_valid,
  input  [2:0]   auto_in_3_a_bits_size,
  input  [3:0]   auto_in_3_a_bits_source,
  input  [33:0]  auto_in_3_a_bits_address,
  input  [63:0]  auto_in_3_a_bits_mask,
  input          auto_in_3_d_ready,
  output         auto_in_3_d_valid,
  output [3:0]   auto_in_3_d_bits_source,
  output         auto_in_2_a_ready,
  input          auto_in_2_a_valid,
  input  [2:0]   auto_in_2_a_bits_size,
  input  [3:0]   auto_in_2_a_bits_source,
  input  [33:0]  auto_in_2_a_bits_address,
  input  [63:0]  auto_in_2_a_bits_mask,
  input          auto_in_2_d_ready,
  output         auto_in_2_d_valid,
  output [3:0]   auto_in_2_d_bits_source,
  output         auto_in_1_a_ready,
  input          auto_in_1_a_valid,
  input  [2:0]   auto_in_1_a_bits_size,
  input  [3:0]   auto_in_1_a_bits_source,
  input  [33:0]  auto_in_1_a_bits_address,
  input  [63:0]  auto_in_1_a_bits_mask,
  input          auto_in_1_d_ready,
  output         auto_in_1_d_valid,
  output [3:0]   auto_in_1_d_bits_source,
  output [511:0] auto_in_1_d_bits_data,
  output         auto_in_0_a_ready,
  input          auto_in_0_a_valid,
  input          auto_in_0_a_bits_source,
  input  [33:0]  auto_in_0_a_bits_address,
  input  [63:0]  auto_in_0_a_bits_mask,
  input  [511:0] auto_in_0_a_bits_data,
  input          auto_in_0_d_ready,
  output         auto_in_0_d_valid,
  output         auto_in_0_d_bits_source,
  input          auto_out_a_ready,
  output         auto_out_a_valid,
  output [2:0]   auto_out_a_bits_opcode,
  output [2:0]   auto_out_a_bits_size,
  output [6:0]   auto_out_a_bits_source,
  output [33:0]  auto_out_a_bits_address,
  output [63:0]  auto_out_a_bits_mask,
  output [511:0] auto_out_a_bits_data,
  output         auto_out_d_ready,
  input          auto_out_d_valid,
  input  [6:0]   auto_out_d_bits_source,
  input  [511:0] auto_out_d_bits_data
);
  wire [6:0] _GEN_1 = {{6'd0}, auto_in_0_a_bits_source}; // @[Xbar.scala 240:55]
  wire [6:0] in_0_a_bits_source = _GEN_1 | 7'h40; // @[Xbar.scala 240:55]
  wire [5:0] _GEN_2 = {{2'd0}, auto_in_1_a_bits_source}; // @[Xbar.scala 240:55]
  wire [5:0] _in_1_a_bits_source_T = _GEN_2 | 6'h30; // @[Xbar.scala 240:55]
  wire [5:0] _GEN_3 = {{2'd0}, auto_in_2_a_bits_source}; // @[Xbar.scala 240:55]
  wire [5:0] _in_2_a_bits_source_T = _GEN_3 | 6'h20; // @[Xbar.scala 240:55]
  wire [4:0] _GEN_4 = {{1'd0}, auto_in_3_a_bits_source}; // @[Xbar.scala 240:55]
  wire [4:0] _in_3_a_bits_source_T = _GEN_4 | 5'h10; // @[Xbar.scala 240:55]
  wire  requestDOI_0_0 = auto_out_d_bits_source[6:1] == 6'h20; // @[Parameters.scala 54:32]
  wire  requestDOI_0_1 = auto_out_d_bits_source[6:4] == 3'h3; // @[Parameters.scala 54:32]
  wire  requestDOI_0_2 = auto_out_d_bits_source[6:4] == 3'h2; // @[Parameters.scala 54:32]
  wire  requestDOI_0_3 = auto_out_d_bits_source[6:4] == 3'h1; // @[Parameters.scala 54:32]
  wire  requestDOI_0_4 = auto_out_d_bits_source[6:4] == 3'h0; // @[Parameters.scala 54:32]
  reg  beatsLeft; // @[Arbiter.scala 88:30]
  wire  idle = ~beatsLeft; // @[Arbiter.scala 89:28]
  wire  latch = idle & auto_out_a_ready; // @[Arbiter.scala 90:24]
  wire [4:0] readys_valid = {auto_in_4_a_valid,auto_in_3_a_valid,auto_in_2_a_valid,auto_in_1_a_valid,auto_in_0_a_valid}; // @[Cat.scala 33:92]
  wire  _readys_T_3 = ~reset; // @[Arbiter.scala 23:12]
  reg [4:0] readys_mask; // @[Arbiter.scala 24:23]
  wire [4:0] _readys_filter_T = ~readys_mask; // @[Arbiter.scala 25:30]
  wire [4:0] _readys_filter_T_1 = readys_valid & _readys_filter_T; // @[Arbiter.scala 25:28]
  wire [9:0] readys_filter = {_readys_filter_T_1,auto_in_4_a_valid,auto_in_3_a_valid,auto_in_2_a_valid,auto_in_1_a_valid
    ,auto_in_0_a_valid}; // @[Cat.scala 33:92]
  wire [9:0] _GEN_5 = {{1'd0}, readys_filter[9:1]}; // @[package.scala 254:43]
  wire [9:0] _readys_unready_T_1 = readys_filter | _GEN_5; // @[package.scala 254:43]
  wire [9:0] _GEN_6 = {{2'd0}, _readys_unready_T_1[9:2]}; // @[package.scala 254:43]
  wire [9:0] _readys_unready_T_3 = _readys_unready_T_1 | _GEN_6; // @[package.scala 254:43]
  wire [9:0] _GEN_7 = {{4'd0}, _readys_unready_T_3[9:4]}; // @[package.scala 254:43]
  wire [9:0] _readys_unready_T_5 = _readys_unready_T_3 | _GEN_7; // @[package.scala 254:43]
  wire [9:0] _readys_unready_T_8 = {readys_mask, 5'h0}; // @[Arbiter.scala 26:66]
  wire [9:0] _GEN_8 = {{1'd0}, _readys_unready_T_5[9:1]}; // @[Arbiter.scala 26:58]
  wire [9:0] readys_unready = _GEN_8 | _readys_unready_T_8; // @[Arbiter.scala 26:58]
  wire [4:0] _readys_readys_T_2 = readys_unready[9:5] & readys_unready[4:0]; // @[Arbiter.scala 27:39]
  wire [4:0] readys_readys = ~_readys_readys_T_2; // @[Arbiter.scala 27:18]
  wire [4:0] _readys_mask_T = readys_readys & readys_valid; // @[Arbiter.scala 29:29]
  wire [5:0] _readys_mask_T_1 = {_readys_mask_T, 1'h0}; // @[package.scala 245:48]
  wire [4:0] _readys_mask_T_3 = _readys_mask_T | _readys_mask_T_1[4:0]; // @[package.scala 245:43]
  wire [6:0] _readys_mask_T_4 = {_readys_mask_T_3, 2'h0}; // @[package.scala 245:48]
  wire [4:0] _readys_mask_T_6 = _readys_mask_T_3 | _readys_mask_T_4[4:0]; // @[package.scala 245:43]
  wire [8:0] _readys_mask_T_7 = {_readys_mask_T_6, 4'h0}; // @[package.scala 245:48]
  wire [4:0] _readys_mask_T_9 = _readys_mask_T_6 | _readys_mask_T_7[4:0]; // @[package.scala 245:43]
  wire  readys_0 = readys_readys[0]; // @[Arbiter.scala 96:86]
  wire  readys_1 = readys_readys[1]; // @[Arbiter.scala 96:86]
  wire  readys_2 = readys_readys[2]; // @[Arbiter.scala 96:86]
  wire  readys_3 = readys_readys[3]; // @[Arbiter.scala 96:86]
  wire  readys_4 = readys_readys[4]; // @[Arbiter.scala 96:86]
  wire  earlyWinner_0 = readys_0 & auto_in_0_a_valid; // @[Arbiter.scala 98:79]
  wire  earlyWinner_1 = readys_1 & auto_in_1_a_valid; // @[Arbiter.scala 98:79]
  wire  earlyWinner_2 = readys_2 & auto_in_2_a_valid; // @[Arbiter.scala 98:79]
  wire  earlyWinner_3 = readys_3 & auto_in_3_a_valid; // @[Arbiter.scala 98:79]
  wire  earlyWinner_4 = readys_4 & auto_in_4_a_valid; // @[Arbiter.scala 98:79]
  wire  prefixOR_2 = earlyWinner_0 | earlyWinner_1; // @[Arbiter.scala 105:53]
  wire  prefixOR_3 = prefixOR_2 | earlyWinner_2; // @[Arbiter.scala 105:53]
  wire  prefixOR_4 = prefixOR_3 | earlyWinner_3; // @[Arbiter.scala 105:53]
  wire  _prefixOR_T = prefixOR_4 | earlyWinner_4; // @[Arbiter.scala 105:53]
  wire  _T_25 = auto_in_0_a_valid | auto_in_1_a_valid | auto_in_2_a_valid | auto_in_3_a_valid | auto_in_4_a_valid; // @[Arbiter.scala 108:36]
  wire  _T_26 = ~(auto_in_0_a_valid | auto_in_1_a_valid | auto_in_2_a_valid | auto_in_3_a_valid | auto_in_4_a_valid); // @[Arbiter.scala 108:15]
  reg  state_0; // @[Arbiter.scala 117:26]
  wire  muxStateEarly_0 = idle ? earlyWinner_0 : state_0; // @[Arbiter.scala 118:30]
  reg  state_1; // @[Arbiter.scala 117:26]
  wire  muxStateEarly_1 = idle ? earlyWinner_1 : state_1; // @[Arbiter.scala 118:30]
  reg  state_2; // @[Arbiter.scala 117:26]
  wire  muxStateEarly_2 = idle ? earlyWinner_2 : state_2; // @[Arbiter.scala 118:30]
  reg  state_3; // @[Arbiter.scala 117:26]
  wire  muxStateEarly_3 = idle ? earlyWinner_3 : state_3; // @[Arbiter.scala 118:30]
  reg  state_4; // @[Arbiter.scala 117:26]
  wire  muxStateEarly_4 = idle ? earlyWinner_4 : state_4; // @[Arbiter.scala 118:30]
  wire  _out_0_a_earlyValid_T_12 = state_0 & auto_in_0_a_valid | state_1 & auto_in_1_a_valid | state_2 &
    auto_in_2_a_valid | state_3 & auto_in_3_a_valid | state_4 & auto_in_4_a_valid; // @[Mux.scala 27:73]
  wire  out_5_0_a_earlyValid = idle ? _T_25 : _out_0_a_earlyValid_T_12; // @[Arbiter.scala 126:29]
  wire  _beatsLeft_T_2 = auto_out_a_ready & out_5_0_a_earlyValid; // @[ReadyValidCancel.scala 49:33]
  wire  allowed_0 = idle ? readys_0 : state_0; // @[Arbiter.scala 122:24]
  wire  allowed_1 = idle ? readys_1 : state_1; // @[Arbiter.scala 122:24]
  wire  allowed_2 = idle ? readys_2 : state_2; // @[Arbiter.scala 122:24]
  wire  allowed_3 = idle ? readys_3 : state_3; // @[Arbiter.scala 122:24]
  wire  allowed_4 = idle ? readys_4 : state_4; // @[Arbiter.scala 122:24]
  wire [63:0] _T_66 = muxStateEarly_0 ? auto_in_0_a_bits_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_67 = muxStateEarly_1 ? auto_in_1_a_bits_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_68 = muxStateEarly_2 ? auto_in_2_a_bits_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_69 = muxStateEarly_3 ? auto_in_3_a_bits_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_70 = muxStateEarly_4 ? auto_in_4_a_bits_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_71 = _T_66 | _T_67; // @[Mux.scala 27:73]
  wire [63:0] _T_72 = _T_71 | _T_68; // @[Mux.scala 27:73]
  wire [63:0] _T_73 = _T_72 | _T_69; // @[Mux.scala 27:73]
  wire [33:0] _T_75 = muxStateEarly_0 ? auto_in_0_a_bits_address : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _T_76 = muxStateEarly_1 ? auto_in_1_a_bits_address : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _T_77 = muxStateEarly_2 ? auto_in_2_a_bits_address : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _T_78 = muxStateEarly_3 ? auto_in_3_a_bits_address : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _T_79 = muxStateEarly_4 ? auto_in_4_a_bits_address : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _T_80 = _T_75 | _T_76; // @[Mux.scala 27:73]
  wire [33:0] _T_81 = _T_80 | _T_77; // @[Mux.scala 27:73]
  wire [33:0] _T_82 = _T_81 | _T_78; // @[Mux.scala 27:73]
  wire [6:0] _T_84 = muxStateEarly_0 ? in_0_a_bits_source : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] in_1_a_bits_source = {{1'd0}, _in_1_a_bits_source_T}; // @[Xbar.scala 234:18 240:29]
  wire [6:0] _T_85 = muxStateEarly_1 ? in_1_a_bits_source : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] in_2_a_bits_source = {{1'd0}, _in_2_a_bits_source_T}; // @[Xbar.scala 234:18 240:29]
  wire [6:0] _T_86 = muxStateEarly_2 ? in_2_a_bits_source : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] in_3_a_bits_source = {{2'd0}, _in_3_a_bits_source_T}; // @[Xbar.scala 234:18 240:29]
  wire [6:0] _T_87 = muxStateEarly_3 ? in_3_a_bits_source : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] in_4_a_bits_source = {{3'd0}, auto_in_4_a_bits_source}; // @[Xbar.scala 234:18 240:29]
  wire [6:0] _T_88 = muxStateEarly_4 ? in_4_a_bits_source : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _T_89 = _T_84 | _T_85; // @[Mux.scala 27:73]
  wire [6:0] _T_90 = _T_89 | _T_86; // @[Mux.scala 27:73]
  wire [6:0] _T_91 = _T_90 | _T_87; // @[Mux.scala 27:73]
  wire [2:0] _T_93 = muxStateEarly_0 ? 3'h6 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_94 = muxStateEarly_1 ? auto_in_1_a_bits_size : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_95 = muxStateEarly_2 ? auto_in_2_a_bits_size : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_96 = muxStateEarly_3 ? auto_in_3_a_bits_size : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_97 = muxStateEarly_4 ? auto_in_4_a_bits_size : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_98 = _T_93 | _T_94; // @[Mux.scala 27:73]
  wire [2:0] _T_99 = _T_98 | _T_95; // @[Mux.scala 27:73]
  wire [2:0] _T_100 = _T_99 | _T_96; // @[Mux.scala 27:73]
  wire [2:0] _T_111 = muxStateEarly_0 ? 3'h1 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_112 = muxStateEarly_1 ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_113 = muxStateEarly_2 ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_114 = muxStateEarly_3 ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_115 = muxStateEarly_4 ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_116 = _T_111 | _T_112; // @[Mux.scala 27:73]
  wire [2:0] _T_117 = _T_116 | _T_113; // @[Mux.scala 27:73]
  wire [2:0] _T_118 = _T_117 | _T_114; // @[Mux.scala 27:73]
  assign auto_in_4_a_ready = auto_out_a_ready & allowed_4; // @[Arbiter.scala 124:31]
  assign auto_in_4_d_valid = auto_out_d_valid & requestDOI_0_4; // @[Xbar.scala 182:40]
  assign auto_in_4_d_bits_source = auto_out_d_bits_source[3:0]; // @[Xbar.scala 231:69]
  assign auto_in_3_a_ready = auto_out_a_ready & allowed_3; // @[Arbiter.scala 124:31]
  assign auto_in_3_d_valid = auto_out_d_valid & requestDOI_0_3; // @[Xbar.scala 182:40]
  assign auto_in_3_d_bits_source = auto_out_d_bits_source[3:0]; // @[Xbar.scala 231:69]
  assign auto_in_2_a_ready = auto_out_a_ready & allowed_2; // @[Arbiter.scala 124:31]
  assign auto_in_2_d_valid = auto_out_d_valid & requestDOI_0_2; // @[Xbar.scala 182:40]
  assign auto_in_2_d_bits_source = auto_out_d_bits_source[3:0]; // @[Xbar.scala 231:69]
  assign auto_in_1_a_ready = auto_out_a_ready & allowed_1; // @[Arbiter.scala 124:31]
  assign auto_in_1_d_valid = auto_out_d_valid & requestDOI_0_1; // @[Xbar.scala 182:40]
  assign auto_in_1_d_bits_source = auto_out_d_bits_source[3:0]; // @[Xbar.scala 231:69]
  assign auto_in_1_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_0_a_ready = auto_out_a_ready & allowed_0; // @[Arbiter.scala 124:31]
  assign auto_in_0_d_valid = auto_out_d_valid & requestDOI_0_0; // @[Xbar.scala 182:40]
  assign auto_in_0_d_bits_source = auto_out_d_bits_source[0]; // @[Xbar.scala 231:69]
  assign auto_out_a_valid = idle ? _T_25 : _out_0_a_earlyValid_T_12; // @[Arbiter.scala 126:29]
  assign auto_out_a_bits_opcode = _T_118 | _T_115; // @[Mux.scala 27:73]
  assign auto_out_a_bits_size = _T_100 | _T_97; // @[Mux.scala 27:73]
  assign auto_out_a_bits_source = _T_91 | _T_88; // @[Mux.scala 27:73]
  assign auto_out_a_bits_address = _T_82 | _T_79; // @[Mux.scala 27:73]
  assign auto_out_a_bits_mask = _T_73 | _T_70; // @[Mux.scala 27:73]
  assign auto_out_a_bits_data = muxStateEarly_0 ? auto_in_0_a_bits_data : 512'h0; // @[Mux.scala 27:73]
  assign auto_out_d_ready = requestDOI_0_0 & auto_in_0_d_ready | requestDOI_0_1 & auto_in_1_d_ready | requestDOI_0_2 &
    auto_in_2_d_ready | requestDOI_0_3 & auto_in_3_d_ready | requestDOI_0_4 & auto_in_4_d_ready; // @[Mux.scala 27:73]
  always @(posedge clock) begin
    if (reset) begin // @[Arbiter.scala 88:30]
      beatsLeft <= 1'h0; // @[Arbiter.scala 88:30]
    end else if (latch) begin // @[Arbiter.scala 114:23]
      beatsLeft <= 1'h0;
    end else begin
      beatsLeft <= beatsLeft - _beatsLeft_T_2;
    end
    if (reset) begin // @[Arbiter.scala 24:23]
      readys_mask <= 5'h1f; // @[Arbiter.scala 24:23]
    end else if (latch & |readys_valid) begin // @[Arbiter.scala 28:32]
      readys_mask <= _readys_mask_T_9; // @[Arbiter.scala 29:12]
    end
    if (reset) begin // @[Arbiter.scala 117:26]
      state_0 <= 1'h0; // @[Arbiter.scala 117:26]
    end else if (idle) begin // @[Arbiter.scala 118:30]
      state_0 <= earlyWinner_0;
    end
    if (reset) begin // @[Arbiter.scala 117:26]
      state_1 <= 1'h0; // @[Arbiter.scala 117:26]
    end else if (idle) begin // @[Arbiter.scala 118:30]
      state_1 <= earlyWinner_1;
    end
    if (reset) begin // @[Arbiter.scala 117:26]
      state_2 <= 1'h0; // @[Arbiter.scala 117:26]
    end else if (idle) begin // @[Arbiter.scala 118:30]
      state_2 <= earlyWinner_2;
    end
    if (reset) begin // @[Arbiter.scala 117:26]
      state_3 <= 1'h0; // @[Arbiter.scala 117:26]
    end else if (idle) begin // @[Arbiter.scala 118:30]
      state_3 <= earlyWinner_3;
    end
    if (reset) begin // @[Arbiter.scala 117:26]
      state_4 <= 1'h0; // @[Arbiter.scala 117:26]
    end else if (idle) begin // @[Arbiter.scala 118:30]
      state_4 <= earlyWinner_4;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_readys_T_3 & ~((~earlyWinner_0 | ~earlyWinner_1) & (~prefixOR_2 | ~earlyWinner_2) & (~prefixOR_3 | ~
          earlyWinner_3) & (~prefixOR_4 | ~earlyWinner_4))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:106 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[Arbiter.scala 106:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~((~earlyWinner_0 | ~earlyWinner_1) & (~prefixOR_2 | ~earlyWinner_2) & (~prefixOR_3 | ~earlyWinner_3) & (~
          prefixOR_4 | ~earlyWinner_4)) & _readys_T_3) begin
          $fatal; // @[Arbiter.scala 106:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_readys_T_3 & ~(~(auto_in_0_a_valid | auto_in_1_a_valid | auto_in_2_a_valid | auto_in_3_a_valid |
          auto_in_4_a_valid) | _prefixOR_T)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:108 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"
            ); // @[Arbiter.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(auto_in_0_a_valid | auto_in_1_a_valid | auto_in_2_a_valid | auto_in_3_a_valid | auto_in_4_a_valid) |
          _prefixOR_T) & _readys_T_3) begin
          $fatal; // @[Arbiter.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_readys_T_3 & ~(_T_26 | _T_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:109 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"
            ); // @[Arbiter.scala 109:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_26 | _T_25) & _readys_T_3) begin
          $fatal; // @[Arbiter.scala 109:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComposerAccSystem(
  input          clock,
  input          reset,
  input          auto_mem_out_a_ready,
  output         auto_mem_out_a_valid,
  output [2:0]   auto_mem_out_a_bits_opcode,
  output [2:0]   auto_mem_out_a_bits_size,
  output [6:0]   auto_mem_out_a_bits_source,
  output [33:0]  auto_mem_out_a_bits_address,
  output [63:0]  auto_mem_out_a_bits_mask,
  output [511:0] auto_mem_out_a_bits_data,
  output         auto_mem_out_d_ready,
  input          auto_mem_out_d_valid,
  input  [6:0]   auto_mem_out_d_bits_source,
  input  [511:0] auto_mem_out_d_bits_data,
  output         io_cmd_ready,
  input          io_cmd_valid,
  input  [6:0]   io_cmd_bits_inst_funct,
  input  [4:0]   io_cmd_bits_inst_rs2,
  input  [4:0]   io_cmd_bits_inst_rs1,
  input  [6:0]   io_cmd_bits_inst_opcode,
  input  [63:0]  io_cmd_bits_rs1,
  input  [63:0]  io_cmd_bits_rs2,
  input          io_resp_ready,
  output         io_resp_valid,
  output [4:0]   io_resp_bits_rd,
  output [63:0]  io_resp_bits_data
);
  wire  acc_clock; // @[Accelerator.scala 145:23]
  wire  acc_reset; // @[Accelerator.scala 145:23]
  wire  acc_auto_EnergyCalc_memory_endpoint_identity_out_4_a_ready; // @[Accelerator.scala 145:23]
  wire  acc_auto_EnergyCalc_memory_endpoint_identity_out_4_a_valid; // @[Accelerator.scala 145:23]
  wire [2:0] acc_auto_EnergyCalc_memory_endpoint_identity_out_4_a_bits_size; // @[Accelerator.scala 145:23]
  wire [3:0] acc_auto_EnergyCalc_memory_endpoint_identity_out_4_a_bits_source; // @[Accelerator.scala 145:23]
  wire [33:0] acc_auto_EnergyCalc_memory_endpoint_identity_out_4_a_bits_address; // @[Accelerator.scala 145:23]
  wire [63:0] acc_auto_EnergyCalc_memory_endpoint_identity_out_4_a_bits_mask; // @[Accelerator.scala 145:23]
  wire  acc_auto_EnergyCalc_memory_endpoint_identity_out_4_d_ready; // @[Accelerator.scala 145:23]
  wire  acc_auto_EnergyCalc_memory_endpoint_identity_out_4_d_valid; // @[Accelerator.scala 145:23]
  wire [3:0] acc_auto_EnergyCalc_memory_endpoint_identity_out_4_d_bits_source; // @[Accelerator.scala 145:23]
  wire  acc_auto_EnergyCalc_memory_endpoint_identity_out_3_a_ready; // @[Accelerator.scala 145:23]
  wire  acc_auto_EnergyCalc_memory_endpoint_identity_out_3_a_valid; // @[Accelerator.scala 145:23]
  wire [2:0] acc_auto_EnergyCalc_memory_endpoint_identity_out_3_a_bits_size; // @[Accelerator.scala 145:23]
  wire [3:0] acc_auto_EnergyCalc_memory_endpoint_identity_out_3_a_bits_source; // @[Accelerator.scala 145:23]
  wire [33:0] acc_auto_EnergyCalc_memory_endpoint_identity_out_3_a_bits_address; // @[Accelerator.scala 145:23]
  wire [63:0] acc_auto_EnergyCalc_memory_endpoint_identity_out_3_a_bits_mask; // @[Accelerator.scala 145:23]
  wire  acc_auto_EnergyCalc_memory_endpoint_identity_out_3_d_ready; // @[Accelerator.scala 145:23]
  wire  acc_auto_EnergyCalc_memory_endpoint_identity_out_3_d_valid; // @[Accelerator.scala 145:23]
  wire [3:0] acc_auto_EnergyCalc_memory_endpoint_identity_out_3_d_bits_source; // @[Accelerator.scala 145:23]
  wire  acc_auto_EnergyCalc_memory_endpoint_identity_out_2_a_ready; // @[Accelerator.scala 145:23]
  wire  acc_auto_EnergyCalc_memory_endpoint_identity_out_2_a_valid; // @[Accelerator.scala 145:23]
  wire [2:0] acc_auto_EnergyCalc_memory_endpoint_identity_out_2_a_bits_size; // @[Accelerator.scala 145:23]
  wire [3:0] acc_auto_EnergyCalc_memory_endpoint_identity_out_2_a_bits_source; // @[Accelerator.scala 145:23]
  wire [33:0] acc_auto_EnergyCalc_memory_endpoint_identity_out_2_a_bits_address; // @[Accelerator.scala 145:23]
  wire [63:0] acc_auto_EnergyCalc_memory_endpoint_identity_out_2_a_bits_mask; // @[Accelerator.scala 145:23]
  wire  acc_auto_EnergyCalc_memory_endpoint_identity_out_2_d_ready; // @[Accelerator.scala 145:23]
  wire  acc_auto_EnergyCalc_memory_endpoint_identity_out_2_d_valid; // @[Accelerator.scala 145:23]
  wire [3:0] acc_auto_EnergyCalc_memory_endpoint_identity_out_2_d_bits_source; // @[Accelerator.scala 145:23]
  wire  acc_auto_EnergyCalc_memory_endpoint_identity_out_1_a_ready; // @[Accelerator.scala 145:23]
  wire  acc_auto_EnergyCalc_memory_endpoint_identity_out_1_a_valid; // @[Accelerator.scala 145:23]
  wire [2:0] acc_auto_EnergyCalc_memory_endpoint_identity_out_1_a_bits_size; // @[Accelerator.scala 145:23]
  wire [3:0] acc_auto_EnergyCalc_memory_endpoint_identity_out_1_a_bits_source; // @[Accelerator.scala 145:23]
  wire [33:0] acc_auto_EnergyCalc_memory_endpoint_identity_out_1_a_bits_address; // @[Accelerator.scala 145:23]
  wire [63:0] acc_auto_EnergyCalc_memory_endpoint_identity_out_1_a_bits_mask; // @[Accelerator.scala 145:23]
  wire  acc_auto_EnergyCalc_memory_endpoint_identity_out_1_d_ready; // @[Accelerator.scala 145:23]
  wire  acc_auto_EnergyCalc_memory_endpoint_identity_out_1_d_valid; // @[Accelerator.scala 145:23]
  wire [3:0] acc_auto_EnergyCalc_memory_endpoint_identity_out_1_d_bits_source; // @[Accelerator.scala 145:23]
  wire [511:0] acc_auto_EnergyCalc_memory_endpoint_identity_out_1_d_bits_data; // @[Accelerator.scala 145:23]
  wire  acc_auto_EnergyCalc_memory_endpoint_identity_out_0_a_ready; // @[Accelerator.scala 145:23]
  wire  acc_auto_EnergyCalc_memory_endpoint_identity_out_0_a_valid; // @[Accelerator.scala 145:23]
  wire  acc_auto_EnergyCalc_memory_endpoint_identity_out_0_a_bits_source; // @[Accelerator.scala 145:23]
  wire [33:0] acc_auto_EnergyCalc_memory_endpoint_identity_out_0_a_bits_address; // @[Accelerator.scala 145:23]
  wire [63:0] acc_auto_EnergyCalc_memory_endpoint_identity_out_0_a_bits_mask; // @[Accelerator.scala 145:23]
  wire [511:0] acc_auto_EnergyCalc_memory_endpoint_identity_out_0_a_bits_data; // @[Accelerator.scala 145:23]
  wire  acc_auto_EnergyCalc_memory_endpoint_identity_out_0_d_ready; // @[Accelerator.scala 145:23]
  wire  acc_auto_EnergyCalc_memory_endpoint_identity_out_0_d_valid; // @[Accelerator.scala 145:23]
  wire  acc_auto_EnergyCalc_memory_endpoint_identity_out_0_d_bits_source; // @[Accelerator.scala 145:23]
  wire  acc_io_cmd_ready; // @[Accelerator.scala 145:23]
  wire  acc_io_cmd_valid; // @[Accelerator.scala 145:23]
  wire [6:0] acc_io_cmd_bits_inst_funct; // @[Accelerator.scala 145:23]
  wire [4:0] acc_io_cmd_bits_inst_rs2; // @[Accelerator.scala 145:23]
  wire [4:0] acc_io_cmd_bits_inst_rs1; // @[Accelerator.scala 145:23]
  wire [6:0] acc_io_cmd_bits_inst_opcode; // @[Accelerator.scala 145:23]
  wire [63:0] acc_io_cmd_bits_rs1; // @[Accelerator.scala 145:23]
  wire [63:0] acc_io_cmd_bits_rs2; // @[Accelerator.scala 145:23]
  wire  acc_io_resp_ready; // @[Accelerator.scala 145:23]
  wire  acc_io_resp_valid; // @[Accelerator.scala 145:23]
  wire [4:0] acc_io_resp_bits_rd; // @[Accelerator.scala 145:23]
  wire [63:0] acc_io_resp_bits_data; // @[Accelerator.scala 145:23]
  wire  crossbarModule_clock; // @[Accelerator.scala 147:34]
  wire  crossbarModule_reset; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_in_4_a_ready; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_in_4_a_valid; // @[Accelerator.scala 147:34]
  wire [2:0] crossbarModule_auto_in_4_a_bits_size; // @[Accelerator.scala 147:34]
  wire [3:0] crossbarModule_auto_in_4_a_bits_source; // @[Accelerator.scala 147:34]
  wire [33:0] crossbarModule_auto_in_4_a_bits_address; // @[Accelerator.scala 147:34]
  wire [63:0] crossbarModule_auto_in_4_a_bits_mask; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_in_4_d_ready; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_in_4_d_valid; // @[Accelerator.scala 147:34]
  wire [3:0] crossbarModule_auto_in_4_d_bits_source; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_in_3_a_ready; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_in_3_a_valid; // @[Accelerator.scala 147:34]
  wire [2:0] crossbarModule_auto_in_3_a_bits_size; // @[Accelerator.scala 147:34]
  wire [3:0] crossbarModule_auto_in_3_a_bits_source; // @[Accelerator.scala 147:34]
  wire [33:0] crossbarModule_auto_in_3_a_bits_address; // @[Accelerator.scala 147:34]
  wire [63:0] crossbarModule_auto_in_3_a_bits_mask; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_in_3_d_ready; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_in_3_d_valid; // @[Accelerator.scala 147:34]
  wire [3:0] crossbarModule_auto_in_3_d_bits_source; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_in_2_a_ready; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_in_2_a_valid; // @[Accelerator.scala 147:34]
  wire [2:0] crossbarModule_auto_in_2_a_bits_size; // @[Accelerator.scala 147:34]
  wire [3:0] crossbarModule_auto_in_2_a_bits_source; // @[Accelerator.scala 147:34]
  wire [33:0] crossbarModule_auto_in_2_a_bits_address; // @[Accelerator.scala 147:34]
  wire [63:0] crossbarModule_auto_in_2_a_bits_mask; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_in_2_d_ready; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_in_2_d_valid; // @[Accelerator.scala 147:34]
  wire [3:0] crossbarModule_auto_in_2_d_bits_source; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_in_1_a_ready; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_in_1_a_valid; // @[Accelerator.scala 147:34]
  wire [2:0] crossbarModule_auto_in_1_a_bits_size; // @[Accelerator.scala 147:34]
  wire [3:0] crossbarModule_auto_in_1_a_bits_source; // @[Accelerator.scala 147:34]
  wire [33:0] crossbarModule_auto_in_1_a_bits_address; // @[Accelerator.scala 147:34]
  wire [63:0] crossbarModule_auto_in_1_a_bits_mask; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_in_1_d_ready; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_in_1_d_valid; // @[Accelerator.scala 147:34]
  wire [3:0] crossbarModule_auto_in_1_d_bits_source; // @[Accelerator.scala 147:34]
  wire [511:0] crossbarModule_auto_in_1_d_bits_data; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_in_0_a_ready; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_in_0_a_valid; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_in_0_a_bits_source; // @[Accelerator.scala 147:34]
  wire [33:0] crossbarModule_auto_in_0_a_bits_address; // @[Accelerator.scala 147:34]
  wire [63:0] crossbarModule_auto_in_0_a_bits_mask; // @[Accelerator.scala 147:34]
  wire [511:0] crossbarModule_auto_in_0_a_bits_data; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_in_0_d_ready; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_in_0_d_valid; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_in_0_d_bits_source; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_out_a_ready; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_out_a_valid; // @[Accelerator.scala 147:34]
  wire [2:0] crossbarModule_auto_out_a_bits_opcode; // @[Accelerator.scala 147:34]
  wire [2:0] crossbarModule_auto_out_a_bits_size; // @[Accelerator.scala 147:34]
  wire [6:0] crossbarModule_auto_out_a_bits_source; // @[Accelerator.scala 147:34]
  wire [33:0] crossbarModule_auto_out_a_bits_address; // @[Accelerator.scala 147:34]
  wire [63:0] crossbarModule_auto_out_a_bits_mask; // @[Accelerator.scala 147:34]
  wire [511:0] crossbarModule_auto_out_a_bits_data; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_out_d_ready; // @[Accelerator.scala 147:34]
  wire  crossbarModule_auto_out_d_valid; // @[Accelerator.scala 147:34]
  wire [6:0] crossbarModule_auto_out_d_bits_source; // @[Accelerator.scala 147:34]
  wire [511:0] crossbarModule_auto_out_d_bits_data; // @[Accelerator.scala 147:34]
  ComposerAcc acc ( // @[Accelerator.scala 145:23]
    .clock(acc_clock),
    .reset(acc_reset),
    .auto_EnergyCalc_memory_endpoint_identity_out_4_a_ready(acc_auto_EnergyCalc_memory_endpoint_identity_out_4_a_ready),
    .auto_EnergyCalc_memory_endpoint_identity_out_4_a_valid(acc_auto_EnergyCalc_memory_endpoint_identity_out_4_a_valid),
    .auto_EnergyCalc_memory_endpoint_identity_out_4_a_bits_size(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_4_a_bits_size),
    .auto_EnergyCalc_memory_endpoint_identity_out_4_a_bits_source(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_4_a_bits_source),
    .auto_EnergyCalc_memory_endpoint_identity_out_4_a_bits_address(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_4_a_bits_address),
    .auto_EnergyCalc_memory_endpoint_identity_out_4_a_bits_mask(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_4_a_bits_mask),
    .auto_EnergyCalc_memory_endpoint_identity_out_4_d_ready(acc_auto_EnergyCalc_memory_endpoint_identity_out_4_d_ready),
    .auto_EnergyCalc_memory_endpoint_identity_out_4_d_valid(acc_auto_EnergyCalc_memory_endpoint_identity_out_4_d_valid),
    .auto_EnergyCalc_memory_endpoint_identity_out_4_d_bits_source(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_4_d_bits_source),
    .auto_EnergyCalc_memory_endpoint_identity_out_3_a_ready(acc_auto_EnergyCalc_memory_endpoint_identity_out_3_a_ready),
    .auto_EnergyCalc_memory_endpoint_identity_out_3_a_valid(acc_auto_EnergyCalc_memory_endpoint_identity_out_3_a_valid),
    .auto_EnergyCalc_memory_endpoint_identity_out_3_a_bits_size(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_3_a_bits_size),
    .auto_EnergyCalc_memory_endpoint_identity_out_3_a_bits_source(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_3_a_bits_source),
    .auto_EnergyCalc_memory_endpoint_identity_out_3_a_bits_address(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_3_a_bits_address),
    .auto_EnergyCalc_memory_endpoint_identity_out_3_a_bits_mask(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_3_a_bits_mask),
    .auto_EnergyCalc_memory_endpoint_identity_out_3_d_ready(acc_auto_EnergyCalc_memory_endpoint_identity_out_3_d_ready),
    .auto_EnergyCalc_memory_endpoint_identity_out_3_d_valid(acc_auto_EnergyCalc_memory_endpoint_identity_out_3_d_valid),
    .auto_EnergyCalc_memory_endpoint_identity_out_3_d_bits_source(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_3_d_bits_source),
    .auto_EnergyCalc_memory_endpoint_identity_out_2_a_ready(acc_auto_EnergyCalc_memory_endpoint_identity_out_2_a_ready),
    .auto_EnergyCalc_memory_endpoint_identity_out_2_a_valid(acc_auto_EnergyCalc_memory_endpoint_identity_out_2_a_valid),
    .auto_EnergyCalc_memory_endpoint_identity_out_2_a_bits_size(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_2_a_bits_size),
    .auto_EnergyCalc_memory_endpoint_identity_out_2_a_bits_source(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_2_a_bits_source),
    .auto_EnergyCalc_memory_endpoint_identity_out_2_a_bits_address(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_2_a_bits_address),
    .auto_EnergyCalc_memory_endpoint_identity_out_2_a_bits_mask(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_2_a_bits_mask),
    .auto_EnergyCalc_memory_endpoint_identity_out_2_d_ready(acc_auto_EnergyCalc_memory_endpoint_identity_out_2_d_ready),
    .auto_EnergyCalc_memory_endpoint_identity_out_2_d_valid(acc_auto_EnergyCalc_memory_endpoint_identity_out_2_d_valid),
    .auto_EnergyCalc_memory_endpoint_identity_out_2_d_bits_source(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_2_d_bits_source),
    .auto_EnergyCalc_memory_endpoint_identity_out_1_a_ready(acc_auto_EnergyCalc_memory_endpoint_identity_out_1_a_ready),
    .auto_EnergyCalc_memory_endpoint_identity_out_1_a_valid(acc_auto_EnergyCalc_memory_endpoint_identity_out_1_a_valid),
    .auto_EnergyCalc_memory_endpoint_identity_out_1_a_bits_size(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_1_a_bits_size),
    .auto_EnergyCalc_memory_endpoint_identity_out_1_a_bits_source(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_1_a_bits_source),
    .auto_EnergyCalc_memory_endpoint_identity_out_1_a_bits_address(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_1_a_bits_address),
    .auto_EnergyCalc_memory_endpoint_identity_out_1_a_bits_mask(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_1_a_bits_mask),
    .auto_EnergyCalc_memory_endpoint_identity_out_1_d_ready(acc_auto_EnergyCalc_memory_endpoint_identity_out_1_d_ready),
    .auto_EnergyCalc_memory_endpoint_identity_out_1_d_valid(acc_auto_EnergyCalc_memory_endpoint_identity_out_1_d_valid),
    .auto_EnergyCalc_memory_endpoint_identity_out_1_d_bits_source(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_1_d_bits_source),
    .auto_EnergyCalc_memory_endpoint_identity_out_1_d_bits_data(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_1_d_bits_data),
    .auto_EnergyCalc_memory_endpoint_identity_out_0_a_ready(acc_auto_EnergyCalc_memory_endpoint_identity_out_0_a_ready),
    .auto_EnergyCalc_memory_endpoint_identity_out_0_a_valid(acc_auto_EnergyCalc_memory_endpoint_identity_out_0_a_valid),
    .auto_EnergyCalc_memory_endpoint_identity_out_0_a_bits_source(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_0_a_bits_source),
    .auto_EnergyCalc_memory_endpoint_identity_out_0_a_bits_address(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_0_a_bits_address),
    .auto_EnergyCalc_memory_endpoint_identity_out_0_a_bits_mask(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_0_a_bits_mask),
    .auto_EnergyCalc_memory_endpoint_identity_out_0_a_bits_data(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_0_a_bits_data),
    .auto_EnergyCalc_memory_endpoint_identity_out_0_d_ready(acc_auto_EnergyCalc_memory_endpoint_identity_out_0_d_ready),
    .auto_EnergyCalc_memory_endpoint_identity_out_0_d_valid(acc_auto_EnergyCalc_memory_endpoint_identity_out_0_d_valid),
    .auto_EnergyCalc_memory_endpoint_identity_out_0_d_bits_source(
      acc_auto_EnergyCalc_memory_endpoint_identity_out_0_d_bits_source),
    .io_cmd_ready(acc_io_cmd_ready),
    .io_cmd_valid(acc_io_cmd_valid),
    .io_cmd_bits_inst_funct(acc_io_cmd_bits_inst_funct),
    .io_cmd_bits_inst_rs2(acc_io_cmd_bits_inst_rs2),
    .io_cmd_bits_inst_rs1(acc_io_cmd_bits_inst_rs1),
    .io_cmd_bits_inst_opcode(acc_io_cmd_bits_inst_opcode),
    .io_cmd_bits_rs1(acc_io_cmd_bits_rs1),
    .io_cmd_bits_rs2(acc_io_cmd_bits_rs2),
    .io_resp_ready(acc_io_resp_ready),
    .io_resp_valid(acc_io_resp_valid),
    .io_resp_bits_rd(acc_io_resp_bits_rd),
    .io_resp_bits_data(acc_io_resp_bits_data)
  );
  TLXbar crossbarModule ( // @[Accelerator.scala 147:34]
    .clock(crossbarModule_clock),
    .reset(crossbarModule_reset),
    .auto_in_4_a_ready(crossbarModule_auto_in_4_a_ready),
    .auto_in_4_a_valid(crossbarModule_auto_in_4_a_valid),
    .auto_in_4_a_bits_size(crossbarModule_auto_in_4_a_bits_size),
    .auto_in_4_a_bits_source(crossbarModule_auto_in_4_a_bits_source),
    .auto_in_4_a_bits_address(crossbarModule_auto_in_4_a_bits_address),
    .auto_in_4_a_bits_mask(crossbarModule_auto_in_4_a_bits_mask),
    .auto_in_4_d_ready(crossbarModule_auto_in_4_d_ready),
    .auto_in_4_d_valid(crossbarModule_auto_in_4_d_valid),
    .auto_in_4_d_bits_source(crossbarModule_auto_in_4_d_bits_source),
    .auto_in_3_a_ready(crossbarModule_auto_in_3_a_ready),
    .auto_in_3_a_valid(crossbarModule_auto_in_3_a_valid),
    .auto_in_3_a_bits_size(crossbarModule_auto_in_3_a_bits_size),
    .auto_in_3_a_bits_source(crossbarModule_auto_in_3_a_bits_source),
    .auto_in_3_a_bits_address(crossbarModule_auto_in_3_a_bits_address),
    .auto_in_3_a_bits_mask(crossbarModule_auto_in_3_a_bits_mask),
    .auto_in_3_d_ready(crossbarModule_auto_in_3_d_ready),
    .auto_in_3_d_valid(crossbarModule_auto_in_3_d_valid),
    .auto_in_3_d_bits_source(crossbarModule_auto_in_3_d_bits_source),
    .auto_in_2_a_ready(crossbarModule_auto_in_2_a_ready),
    .auto_in_2_a_valid(crossbarModule_auto_in_2_a_valid),
    .auto_in_2_a_bits_size(crossbarModule_auto_in_2_a_bits_size),
    .auto_in_2_a_bits_source(crossbarModule_auto_in_2_a_bits_source),
    .auto_in_2_a_bits_address(crossbarModule_auto_in_2_a_bits_address),
    .auto_in_2_a_bits_mask(crossbarModule_auto_in_2_a_bits_mask),
    .auto_in_2_d_ready(crossbarModule_auto_in_2_d_ready),
    .auto_in_2_d_valid(crossbarModule_auto_in_2_d_valid),
    .auto_in_2_d_bits_source(crossbarModule_auto_in_2_d_bits_source),
    .auto_in_1_a_ready(crossbarModule_auto_in_1_a_ready),
    .auto_in_1_a_valid(crossbarModule_auto_in_1_a_valid),
    .auto_in_1_a_bits_size(crossbarModule_auto_in_1_a_bits_size),
    .auto_in_1_a_bits_source(crossbarModule_auto_in_1_a_bits_source),
    .auto_in_1_a_bits_address(crossbarModule_auto_in_1_a_bits_address),
    .auto_in_1_a_bits_mask(crossbarModule_auto_in_1_a_bits_mask),
    .auto_in_1_d_ready(crossbarModule_auto_in_1_d_ready),
    .auto_in_1_d_valid(crossbarModule_auto_in_1_d_valid),
    .auto_in_1_d_bits_source(crossbarModule_auto_in_1_d_bits_source),
    .auto_in_1_d_bits_data(crossbarModule_auto_in_1_d_bits_data),
    .auto_in_0_a_ready(crossbarModule_auto_in_0_a_ready),
    .auto_in_0_a_valid(crossbarModule_auto_in_0_a_valid),
    .auto_in_0_a_bits_source(crossbarModule_auto_in_0_a_bits_source),
    .auto_in_0_a_bits_address(crossbarModule_auto_in_0_a_bits_address),
    .auto_in_0_a_bits_mask(crossbarModule_auto_in_0_a_bits_mask),
    .auto_in_0_a_bits_data(crossbarModule_auto_in_0_a_bits_data),
    .auto_in_0_d_ready(crossbarModule_auto_in_0_d_ready),
    .auto_in_0_d_valid(crossbarModule_auto_in_0_d_valid),
    .auto_in_0_d_bits_source(crossbarModule_auto_in_0_d_bits_source),
    .auto_out_a_ready(crossbarModule_auto_out_a_ready),
    .auto_out_a_valid(crossbarModule_auto_out_a_valid),
    .auto_out_a_bits_opcode(crossbarModule_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(crossbarModule_auto_out_a_bits_size),
    .auto_out_a_bits_source(crossbarModule_auto_out_a_bits_source),
    .auto_out_a_bits_address(crossbarModule_auto_out_a_bits_address),
    .auto_out_a_bits_mask(crossbarModule_auto_out_a_bits_mask),
    .auto_out_a_bits_data(crossbarModule_auto_out_a_bits_data),
    .auto_out_d_ready(crossbarModule_auto_out_d_ready),
    .auto_out_d_valid(crossbarModule_auto_out_d_valid),
    .auto_out_d_bits_source(crossbarModule_auto_out_d_bits_source),
    .auto_out_d_bits_data(crossbarModule_auto_out_d_bits_data)
  );
  assign auto_mem_out_a_valid = crossbarModule_auto_out_a_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_mem_out_a_bits_opcode = crossbarModule_auto_out_a_bits_opcode; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_mem_out_a_bits_size = crossbarModule_auto_out_a_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_mem_out_a_bits_source = crossbarModule_auto_out_a_bits_source; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_mem_out_a_bits_address = crossbarModule_auto_out_a_bits_address; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_mem_out_a_bits_mask = crossbarModule_auto_out_a_bits_mask; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_mem_out_a_bits_data = crossbarModule_auto_out_a_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_mem_out_d_ready = crossbarModule_auto_out_d_ready; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_cmd_ready = acc_io_cmd_ready; // @[Accelerator.scala 164:27]
  assign io_resp_valid = acc_io_resp_valid; // @[Accelerator.scala 165:11]
  assign io_resp_bits_rd = acc_io_resp_bits_rd; // @[Accelerator.scala 165:11]
  assign io_resp_bits_data = acc_io_resp_bits_data; // @[Accelerator.scala 165:11]
  assign acc_clock = clock;
  assign acc_reset = reset;
  assign acc_auto_EnergyCalc_memory_endpoint_identity_out_4_a_ready = crossbarModule_auto_in_4_a_ready; // @[LazyModule.scala 355:16]
  assign acc_auto_EnergyCalc_memory_endpoint_identity_out_4_d_valid = crossbarModule_auto_in_4_d_valid; // @[LazyModule.scala 355:16]
  assign acc_auto_EnergyCalc_memory_endpoint_identity_out_4_d_bits_source = crossbarModule_auto_in_4_d_bits_source; // @[LazyModule.scala 355:16]
  assign acc_auto_EnergyCalc_memory_endpoint_identity_out_3_a_ready = crossbarModule_auto_in_3_a_ready; // @[LazyModule.scala 355:16]
  assign acc_auto_EnergyCalc_memory_endpoint_identity_out_3_d_valid = crossbarModule_auto_in_3_d_valid; // @[LazyModule.scala 355:16]
  assign acc_auto_EnergyCalc_memory_endpoint_identity_out_3_d_bits_source = crossbarModule_auto_in_3_d_bits_source; // @[LazyModule.scala 355:16]
  assign acc_auto_EnergyCalc_memory_endpoint_identity_out_2_a_ready = crossbarModule_auto_in_2_a_ready; // @[LazyModule.scala 355:16]
  assign acc_auto_EnergyCalc_memory_endpoint_identity_out_2_d_valid = crossbarModule_auto_in_2_d_valid; // @[LazyModule.scala 355:16]
  assign acc_auto_EnergyCalc_memory_endpoint_identity_out_2_d_bits_source = crossbarModule_auto_in_2_d_bits_source; // @[LazyModule.scala 355:16]
  assign acc_auto_EnergyCalc_memory_endpoint_identity_out_1_a_ready = crossbarModule_auto_in_1_a_ready; // @[LazyModule.scala 355:16]
  assign acc_auto_EnergyCalc_memory_endpoint_identity_out_1_d_valid = crossbarModule_auto_in_1_d_valid; // @[LazyModule.scala 355:16]
  assign acc_auto_EnergyCalc_memory_endpoint_identity_out_1_d_bits_source = crossbarModule_auto_in_1_d_bits_source; // @[LazyModule.scala 355:16]
  assign acc_auto_EnergyCalc_memory_endpoint_identity_out_1_d_bits_data = crossbarModule_auto_in_1_d_bits_data; // @[LazyModule.scala 355:16]
  assign acc_auto_EnergyCalc_memory_endpoint_identity_out_0_a_ready = crossbarModule_auto_in_0_a_ready; // @[LazyModule.scala 355:16]
  assign acc_auto_EnergyCalc_memory_endpoint_identity_out_0_d_valid = crossbarModule_auto_in_0_d_valid; // @[LazyModule.scala 355:16]
  assign acc_auto_EnergyCalc_memory_endpoint_identity_out_0_d_bits_source = crossbarModule_auto_in_0_d_bits_source; // @[LazyModule.scala 355:16]
  assign acc_io_cmd_valid = io_cmd_valid; // @[Accelerator.scala 164:27]
  assign acc_io_cmd_bits_inst_funct = io_cmd_bits_inst_funct; // @[Accelerator.scala 164:27]
  assign acc_io_cmd_bits_inst_rs2 = io_cmd_bits_inst_rs2; // @[Accelerator.scala 164:27]
  assign acc_io_cmd_bits_inst_rs1 = io_cmd_bits_inst_rs1; // @[Accelerator.scala 164:27]
  assign acc_io_cmd_bits_inst_opcode = io_cmd_bits_inst_opcode; // @[Accelerator.scala 164:27]
  assign acc_io_cmd_bits_rs1 = io_cmd_bits_rs1; // @[Accelerator.scala 164:27]
  assign acc_io_cmd_bits_rs2 = io_cmd_bits_rs2; // @[Accelerator.scala 164:27]
  assign acc_io_resp_ready = io_resp_ready; // @[Accelerator.scala 165:11]
  assign crossbarModule_clock = clock;
  assign crossbarModule_reset = reset;
  assign crossbarModule_auto_in_4_a_valid = acc_auto_EnergyCalc_memory_endpoint_identity_out_4_a_valid; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_4_a_bits_size = acc_auto_EnergyCalc_memory_endpoint_identity_out_4_a_bits_size; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_4_a_bits_source = acc_auto_EnergyCalc_memory_endpoint_identity_out_4_a_bits_source; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_4_a_bits_address = acc_auto_EnergyCalc_memory_endpoint_identity_out_4_a_bits_address; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_4_a_bits_mask = acc_auto_EnergyCalc_memory_endpoint_identity_out_4_a_bits_mask; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_4_d_ready = acc_auto_EnergyCalc_memory_endpoint_identity_out_4_d_ready; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_3_a_valid = acc_auto_EnergyCalc_memory_endpoint_identity_out_3_a_valid; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_3_a_bits_size = acc_auto_EnergyCalc_memory_endpoint_identity_out_3_a_bits_size; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_3_a_bits_source = acc_auto_EnergyCalc_memory_endpoint_identity_out_3_a_bits_source; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_3_a_bits_address = acc_auto_EnergyCalc_memory_endpoint_identity_out_3_a_bits_address; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_3_a_bits_mask = acc_auto_EnergyCalc_memory_endpoint_identity_out_3_a_bits_mask; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_3_d_ready = acc_auto_EnergyCalc_memory_endpoint_identity_out_3_d_ready; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_2_a_valid = acc_auto_EnergyCalc_memory_endpoint_identity_out_2_a_valid; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_2_a_bits_size = acc_auto_EnergyCalc_memory_endpoint_identity_out_2_a_bits_size; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_2_a_bits_source = acc_auto_EnergyCalc_memory_endpoint_identity_out_2_a_bits_source; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_2_a_bits_address = acc_auto_EnergyCalc_memory_endpoint_identity_out_2_a_bits_address; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_2_a_bits_mask = acc_auto_EnergyCalc_memory_endpoint_identity_out_2_a_bits_mask; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_2_d_ready = acc_auto_EnergyCalc_memory_endpoint_identity_out_2_d_ready; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_1_a_valid = acc_auto_EnergyCalc_memory_endpoint_identity_out_1_a_valid; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_1_a_bits_size = acc_auto_EnergyCalc_memory_endpoint_identity_out_1_a_bits_size; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_1_a_bits_source = acc_auto_EnergyCalc_memory_endpoint_identity_out_1_a_bits_source; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_1_a_bits_address = acc_auto_EnergyCalc_memory_endpoint_identity_out_1_a_bits_address; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_1_a_bits_mask = acc_auto_EnergyCalc_memory_endpoint_identity_out_1_a_bits_mask; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_1_d_ready = acc_auto_EnergyCalc_memory_endpoint_identity_out_1_d_ready; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_0_a_valid = acc_auto_EnergyCalc_memory_endpoint_identity_out_0_a_valid; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_0_a_bits_source = acc_auto_EnergyCalc_memory_endpoint_identity_out_0_a_bits_source; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_0_a_bits_address = acc_auto_EnergyCalc_memory_endpoint_identity_out_0_a_bits_address; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_0_a_bits_mask = acc_auto_EnergyCalc_memory_endpoint_identity_out_0_a_bits_mask; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_0_a_bits_data = acc_auto_EnergyCalc_memory_endpoint_identity_out_0_a_bits_data; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_in_0_d_ready = acc_auto_EnergyCalc_memory_endpoint_identity_out_0_d_ready; // @[LazyModule.scala 355:16]
  assign crossbarModule_auto_out_a_ready = auto_mem_out_a_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign crossbarModule_auto_out_d_valid = auto_mem_out_d_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign crossbarModule_auto_out_d_bits_source = auto_mem_out_d_bits_source; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign crossbarModule_auto_out_d_bits_data = auto_mem_out_d_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
endmodule
module Queue_6(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [6:0]  io_enq_bits_id,
  input  [33:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_len,
  input  [2:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_burst,
  input         io_enq_bits_lock,
  input  [3:0]  io_enq_bits_cache,
  input  [2:0]  io_enq_bits_prot,
  input  [3:0]  io_enq_bits_qos,
  input  [6:0]  io_enq_bits_echo_tl_state_source,
  input         io_deq_ready,
  output        io_deq_valid,
  output [6:0]  io_deq_bits_id,
  output [33:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_len,
  output [2:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_burst,
  output        io_deq_bits_lock,
  output [3:0]  io_deq_bits_cache,
  output [2:0]  io_deq_bits_prot,
  output [3:0]  io_deq_bits_qos,
  output [6:0]  io_deq_bits_echo_tl_state_source
);
  reg [6:0] ram_id [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [6:0] ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [6:0] ram_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [33:0] ram_addr [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_addr_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_addr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [33:0] ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [33:0] ram_addr_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_addr_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_addr_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_addr_MPORT_en; // @[Decoupled.scala 273:95]
  reg [7:0] ram_len [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_len_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_len_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [7:0] ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [7:0] ram_len_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_len_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_len_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_len_MPORT_en; // @[Decoupled.scala 273:95]
  reg [2:0] ram_size [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_size_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_burst [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_burst_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_burst_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_burst_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_burst_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_burst_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_burst_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_lock [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_lock_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_lock_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_lock_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_lock_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_lock_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_lock_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_lock_MPORT_en; // @[Decoupled.scala 273:95]
  reg [3:0] ram_cache [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_cache_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_cache_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [3:0] ram_cache_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [3:0] ram_cache_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_cache_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_cache_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_cache_MPORT_en; // @[Decoupled.scala 273:95]
  reg [2:0] ram_prot [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_prot_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_prot_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [2:0] ram_prot_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_prot_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_prot_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_prot_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_prot_MPORT_en; // @[Decoupled.scala 273:95]
  reg [3:0] ram_qos [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_qos_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_qos_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [3:0] ram_qos_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [3:0] ram_qos_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_qos_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_qos_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_qos_MPORT_en; // @[Decoupled.scala 273:95]
  reg [6:0] ram_echo_tl_state_source [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [6:0] ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [6:0] ram_echo_tl_state_source_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = enq_ptr_value;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_addr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_addr_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = enq_ptr_value;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_len_io_deq_bits_MPORT_en = 1'h1;
  assign ram_len_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_len_io_deq_bits_MPORT_data = ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_len_MPORT_data = io_enq_bits_len;
  assign ram_len_MPORT_addr = enq_ptr_value;
  assign ram_len_MPORT_mask = 1'h1;
  assign ram_len_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = enq_ptr_value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_burst_io_deq_bits_MPORT_en = 1'h1;
  assign ram_burst_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_burst_io_deq_bits_MPORT_data = ram_burst[ram_burst_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_burst_MPORT_data = io_enq_bits_burst;
  assign ram_burst_MPORT_addr = enq_ptr_value;
  assign ram_burst_MPORT_mask = 1'h1;
  assign ram_burst_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_lock_io_deq_bits_MPORT_en = 1'h1;
  assign ram_lock_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_lock_io_deq_bits_MPORT_data = ram_lock[ram_lock_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_lock_MPORT_data = io_enq_bits_lock;
  assign ram_lock_MPORT_addr = enq_ptr_value;
  assign ram_lock_MPORT_mask = 1'h1;
  assign ram_lock_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_cache_io_deq_bits_MPORT_en = 1'h1;
  assign ram_cache_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_cache_io_deq_bits_MPORT_data = ram_cache[ram_cache_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_cache_MPORT_data = io_enq_bits_cache;
  assign ram_cache_MPORT_addr = enq_ptr_value;
  assign ram_cache_MPORT_mask = 1'h1;
  assign ram_cache_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_prot_io_deq_bits_MPORT_en = 1'h1;
  assign ram_prot_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_prot_io_deq_bits_MPORT_data = ram_prot[ram_prot_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_prot_MPORT_data = io_enq_bits_prot;
  assign ram_prot_MPORT_addr = enq_ptr_value;
  assign ram_prot_MPORT_mask = 1'h1;
  assign ram_prot_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_qos_io_deq_bits_MPORT_en = 1'h1;
  assign ram_qos_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_qos_io_deq_bits_MPORT_data = ram_qos[ram_qos_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_qos_MPORT_data = io_enq_bits_qos;
  assign ram_qos_MPORT_addr = enq_ptr_value;
  assign ram_qos_MPORT_mask = 1'h1;
  assign ram_qos_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_data =
    ram_echo_tl_state_source[ram_echo_tl_state_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_echo_tl_state_source_MPORT_data = io_enq_bits_echo_tl_state_source;
  assign ram_echo_tl_state_source_MPORT_addr = enq_ptr_value;
  assign ram_echo_tl_state_source_MPORT_mask = 1'h1;
  assign ram_echo_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_id = ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_addr = ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_len = ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_burst = ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_lock = ram_lock_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_cache = ram_cache_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_prot = ram_prot_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_qos = ram_qos_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_echo_tl_state_source = ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_len_MPORT_en & ram_len_MPORT_mask) begin
      ram_len[ram_len_MPORT_addr] <= ram_len_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_burst_MPORT_en & ram_burst_MPORT_mask) begin
      ram_burst[ram_burst_MPORT_addr] <= ram_burst_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_lock_MPORT_en & ram_lock_MPORT_mask) begin
      ram_lock[ram_lock_MPORT_addr] <= ram_lock_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_cache_MPORT_en & ram_cache_MPORT_mask) begin
      ram_cache[ram_cache_MPORT_addr] <= ram_cache_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_prot_MPORT_en & ram_prot_MPORT_mask) begin
      ram_prot[ram_prot_MPORT_addr] <= ram_prot_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_qos_MPORT_en & ram_qos_MPORT_mask) begin
      ram_qos[ram_qos_MPORT_addr] <= ram_qos_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_echo_tl_state_source_MPORT_en & ram_echo_tl_state_source_MPORT_mask) begin
      ram_echo_tl_state_source[ram_echo_tl_state_source_MPORT_addr] <= ram_echo_tl_state_source_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
endmodule
module Queue_7(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [511:0] io_enq_bits_data,
  input  [63:0]  io_enq_bits_strb,
  input          io_enq_bits_last,
  input          io_deq_ready,
  output         io_deq_valid,
  output [511:0] io_deq_bits_data,
  output [63:0]  io_deq_bits_strb,
  output         io_deq_bits_last
);
  reg [511:0] ram_data [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [511:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [511:0] ram_data_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 273:95]
  reg [63:0] ram_strb [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_strb_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_strb_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [63:0] ram_strb_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [63:0] ram_strb_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_strb_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_strb_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_strb_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_last [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_strb_io_deq_bits_MPORT_en = 1'h1;
  assign ram_strb_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_strb_io_deq_bits_MPORT_data = ram_strb[ram_strb_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_strb_MPORT_data = io_enq_bits_strb;
  assign ram_strb_MPORT_addr = enq_ptr_value;
  assign ram_strb_MPORT_mask = 1'h1;
  assign ram_strb_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_last_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_last_io_deq_bits_MPORT_data = ram_last[ram_last_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_last_MPORT_data = io_enq_bits_last;
  assign ram_last_MPORT_addr = enq_ptr_value;
  assign ram_last_MPORT_mask = 1'h1;
  assign ram_last_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_strb = ram_strb_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_last = ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_strb_MPORT_en & ram_strb_MPORT_mask) begin
      ram_strb[ram_strb_MPORT_addr] <= ram_strb_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_last_MPORT_en & ram_last_MPORT_mask) begin
      ram_last[ram_last_MPORT_addr] <= ram_last_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
endmodule
module Queue_8(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [6:0] io_enq_bits_id,
  input  [6:0] io_enq_bits_echo_tl_state_source,
  input        io_deq_ready,
  output       io_deq_valid,
  output [6:0] io_deq_bits_id,
  output [6:0] io_deq_bits_echo_tl_state_source
);
  reg [6:0] ram_id [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [6:0] ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [6:0] ram_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [6:0] ram_echo_tl_state_source [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [6:0] ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [6:0] ram_echo_tl_state_source_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = enq_ptr_value;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_data =
    ram_echo_tl_state_source[ram_echo_tl_state_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_echo_tl_state_source_MPORT_data = io_enq_bits_echo_tl_state_source;
  assign ram_echo_tl_state_source_MPORT_addr = enq_ptr_value;
  assign ram_echo_tl_state_source_MPORT_mask = 1'h1;
  assign ram_echo_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_id = ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_echo_tl_state_source = ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_echo_tl_state_source_MPORT_en & ram_echo_tl_state_source_MPORT_mask) begin
      ram_echo_tl_state_source[ram_echo_tl_state_source_MPORT_addr] <= ram_echo_tl_state_source_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
endmodule
module Queue_10(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [6:0]   io_enq_bits_id,
  input  [511:0] io_enq_bits_data,
  input  [6:0]   io_enq_bits_echo_tl_state_source,
  input          io_enq_bits_last,
  input          io_deq_ready,
  output         io_deq_valid,
  output [6:0]   io_deq_bits_id,
  output [511:0] io_deq_bits_data,
  output [6:0]   io_deq_bits_echo_tl_state_source,
  output         io_deq_bits_last
);
  reg [6:0] ram_id [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [6:0] ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [6:0] ram_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [511:0] ram_data [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [511:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [511:0] ram_data_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 273:95]
  reg [6:0] ram_echo_tl_state_source [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [6:0] ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [6:0] ram_echo_tl_state_source_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_last [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = enq_ptr_value;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_data =
    ram_echo_tl_state_source[ram_echo_tl_state_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_echo_tl_state_source_MPORT_data = io_enq_bits_echo_tl_state_source;
  assign ram_echo_tl_state_source_MPORT_addr = enq_ptr_value;
  assign ram_echo_tl_state_source_MPORT_mask = 1'h1;
  assign ram_echo_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_last_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_last_io_deq_bits_MPORT_data = ram_last[ram_last_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_last_MPORT_data = io_enq_bits_last;
  assign ram_last_MPORT_addr = enq_ptr_value;
  assign ram_last_MPORT_mask = 1'h1;
  assign ram_last_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_id = ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_echo_tl_state_source = ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_last = ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_echo_tl_state_source_MPORT_en & ram_echo_tl_state_source_MPORT_mask) begin
      ram_echo_tl_state_source[ram_echo_tl_state_source_MPORT_addr] <= ram_echo_tl_state_source_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_last_MPORT_en & ram_last_MPORT_mask) begin
      ram_last[ram_last_MPORT_addr] <= ram_last_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
endmodule
module AXI4Buffer(
  input          clock,
  input          reset,
  output         auto_in_aw_ready,
  input          auto_in_aw_valid,
  input  [6:0]   auto_in_aw_bits_id,
  input  [33:0]  auto_in_aw_bits_addr,
  input  [7:0]   auto_in_aw_bits_len,
  input  [2:0]   auto_in_aw_bits_size,
  input  [1:0]   auto_in_aw_bits_burst,
  input          auto_in_aw_bits_lock,
  input  [3:0]   auto_in_aw_bits_cache,
  input  [2:0]   auto_in_aw_bits_prot,
  input  [3:0]   auto_in_aw_bits_qos,
  input  [6:0]   auto_in_aw_bits_echo_tl_state_source,
  output         auto_in_w_ready,
  input          auto_in_w_valid,
  input  [511:0] auto_in_w_bits_data,
  input  [63:0]  auto_in_w_bits_strb,
  input          auto_in_w_bits_last,
  input          auto_in_b_ready,
  output         auto_in_b_valid,
  output [6:0]   auto_in_b_bits_id,
  output [6:0]   auto_in_b_bits_echo_tl_state_source,
  output         auto_in_ar_ready,
  input          auto_in_ar_valid,
  input  [6:0]   auto_in_ar_bits_id,
  input  [33:0]  auto_in_ar_bits_addr,
  input  [7:0]   auto_in_ar_bits_len,
  input  [2:0]   auto_in_ar_bits_size,
  input  [1:0]   auto_in_ar_bits_burst,
  input          auto_in_ar_bits_lock,
  input  [3:0]   auto_in_ar_bits_cache,
  input  [2:0]   auto_in_ar_bits_prot,
  input  [3:0]   auto_in_ar_bits_qos,
  input  [6:0]   auto_in_ar_bits_echo_tl_state_source,
  input          auto_in_r_ready,
  output         auto_in_r_valid,
  output [6:0]   auto_in_r_bits_id,
  output [511:0] auto_in_r_bits_data,
  output [6:0]   auto_in_r_bits_echo_tl_state_source,
  output         auto_in_r_bits_last,
  input          auto_out_aw_ready,
  output         auto_out_aw_valid,
  output [6:0]   auto_out_aw_bits_id,
  output [33:0]  auto_out_aw_bits_addr,
  output [7:0]   auto_out_aw_bits_len,
  output [2:0]   auto_out_aw_bits_size,
  output [1:0]   auto_out_aw_bits_burst,
  output         auto_out_aw_bits_lock,
  output [3:0]   auto_out_aw_bits_cache,
  output [2:0]   auto_out_aw_bits_prot,
  output [3:0]   auto_out_aw_bits_qos,
  output [6:0]   auto_out_aw_bits_echo_tl_state_source,
  input          auto_out_w_ready,
  output         auto_out_w_valid,
  output [511:0] auto_out_w_bits_data,
  output [63:0]  auto_out_w_bits_strb,
  output         auto_out_w_bits_last,
  output         auto_out_b_ready,
  input          auto_out_b_valid,
  input  [6:0]   auto_out_b_bits_id,
  input  [6:0]   auto_out_b_bits_echo_tl_state_source,
  input          auto_out_ar_ready,
  output         auto_out_ar_valid,
  output [6:0]   auto_out_ar_bits_id,
  output [33:0]  auto_out_ar_bits_addr,
  output [7:0]   auto_out_ar_bits_len,
  output [2:0]   auto_out_ar_bits_size,
  output [1:0]   auto_out_ar_bits_burst,
  output         auto_out_ar_bits_lock,
  output [3:0]   auto_out_ar_bits_cache,
  output [2:0]   auto_out_ar_bits_prot,
  output [3:0]   auto_out_ar_bits_qos,
  output [6:0]   auto_out_ar_bits_echo_tl_state_source,
  output         auto_out_r_ready,
  input          auto_out_r_valid,
  input  [6:0]   auto_out_r_bits_id,
  input  [511:0] auto_out_r_bits_data,
  input  [6:0]   auto_out_r_bits_echo_tl_state_source,
  input          auto_out_r_bits_last
);
  wire  x1_aw_deq_clock; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_reset; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [6:0] x1_aw_deq_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire [33:0] x1_aw_deq_io_enq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] x1_aw_deq_io_enq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] x1_aw_deq_io_enq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] x1_aw_deq_io_enq_bits_burst; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_enq_bits_lock; // @[Decoupled.scala 375:21]
  wire [3:0] x1_aw_deq_io_enq_bits_cache; // @[Decoupled.scala 375:21]
  wire [2:0] x1_aw_deq_io_enq_bits_prot; // @[Decoupled.scala 375:21]
  wire [3:0] x1_aw_deq_io_enq_bits_qos; // @[Decoupled.scala 375:21]
  wire [6:0] x1_aw_deq_io_enq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [6:0] x1_aw_deq_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [33:0] x1_aw_deq_io_deq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] x1_aw_deq_io_deq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] x1_aw_deq_io_deq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] x1_aw_deq_io_deq_bits_burst; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_deq_bits_lock; // @[Decoupled.scala 375:21]
  wire [3:0] x1_aw_deq_io_deq_bits_cache; // @[Decoupled.scala 375:21]
  wire [2:0] x1_aw_deq_io_deq_bits_prot; // @[Decoupled.scala 375:21]
  wire [3:0] x1_aw_deq_io_deq_bits_qos; // @[Decoupled.scala 375:21]
  wire [6:0] x1_aw_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_clock; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_reset; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [511:0] x1_w_deq_io_enq_bits_data; // @[Decoupled.scala 375:21]
  wire [63:0] x1_w_deq_io_enq_bits_strb; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_enq_bits_last; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [511:0] x1_w_deq_io_deq_bits_data; // @[Decoupled.scala 375:21]
  wire [63:0] x1_w_deq_io_deq_bits_strb; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_deq_bits_last; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_clock; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_reset; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [6:0] bundleIn_0_b_deq_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire [6:0] bundleIn_0_b_deq_io_enq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [6:0] bundleIn_0_b_deq_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [6:0] bundleIn_0_b_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_clock; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_reset; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [6:0] x1_ar_deq_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire [33:0] x1_ar_deq_io_enq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] x1_ar_deq_io_enq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] x1_ar_deq_io_enq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] x1_ar_deq_io_enq_bits_burst; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_enq_bits_lock; // @[Decoupled.scala 375:21]
  wire [3:0] x1_ar_deq_io_enq_bits_cache; // @[Decoupled.scala 375:21]
  wire [2:0] x1_ar_deq_io_enq_bits_prot; // @[Decoupled.scala 375:21]
  wire [3:0] x1_ar_deq_io_enq_bits_qos; // @[Decoupled.scala 375:21]
  wire [6:0] x1_ar_deq_io_enq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [6:0] x1_ar_deq_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [33:0] x1_ar_deq_io_deq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] x1_ar_deq_io_deq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] x1_ar_deq_io_deq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] x1_ar_deq_io_deq_bits_burst; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_deq_bits_lock; // @[Decoupled.scala 375:21]
  wire [3:0] x1_ar_deq_io_deq_bits_cache; // @[Decoupled.scala 375:21]
  wire [2:0] x1_ar_deq_io_deq_bits_prot; // @[Decoupled.scala 375:21]
  wire [3:0] x1_ar_deq_io_deq_bits_qos; // @[Decoupled.scala 375:21]
  wire [6:0] x1_ar_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_clock; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_reset; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [6:0] bundleIn_0_r_deq_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire [511:0] bundleIn_0_r_deq_io_enq_bits_data; // @[Decoupled.scala 375:21]
  wire [6:0] bundleIn_0_r_deq_io_enq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_enq_bits_last; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [6:0] bundleIn_0_r_deq_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [511:0] bundleIn_0_r_deq_io_deq_bits_data; // @[Decoupled.scala 375:21]
  wire [6:0] bundleIn_0_r_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_deq_bits_last; // @[Decoupled.scala 375:21]
  Queue_6 x1_aw_deq ( // @[Decoupled.scala 375:21]
    .clock(x1_aw_deq_clock),
    .reset(x1_aw_deq_reset),
    .io_enq_ready(x1_aw_deq_io_enq_ready),
    .io_enq_valid(x1_aw_deq_io_enq_valid),
    .io_enq_bits_id(x1_aw_deq_io_enq_bits_id),
    .io_enq_bits_addr(x1_aw_deq_io_enq_bits_addr),
    .io_enq_bits_len(x1_aw_deq_io_enq_bits_len),
    .io_enq_bits_size(x1_aw_deq_io_enq_bits_size),
    .io_enq_bits_burst(x1_aw_deq_io_enq_bits_burst),
    .io_enq_bits_lock(x1_aw_deq_io_enq_bits_lock),
    .io_enq_bits_cache(x1_aw_deq_io_enq_bits_cache),
    .io_enq_bits_prot(x1_aw_deq_io_enq_bits_prot),
    .io_enq_bits_qos(x1_aw_deq_io_enq_bits_qos),
    .io_enq_bits_echo_tl_state_source(x1_aw_deq_io_enq_bits_echo_tl_state_source),
    .io_deq_ready(x1_aw_deq_io_deq_ready),
    .io_deq_valid(x1_aw_deq_io_deq_valid),
    .io_deq_bits_id(x1_aw_deq_io_deq_bits_id),
    .io_deq_bits_addr(x1_aw_deq_io_deq_bits_addr),
    .io_deq_bits_len(x1_aw_deq_io_deq_bits_len),
    .io_deq_bits_size(x1_aw_deq_io_deq_bits_size),
    .io_deq_bits_burst(x1_aw_deq_io_deq_bits_burst),
    .io_deq_bits_lock(x1_aw_deq_io_deq_bits_lock),
    .io_deq_bits_cache(x1_aw_deq_io_deq_bits_cache),
    .io_deq_bits_prot(x1_aw_deq_io_deq_bits_prot),
    .io_deq_bits_qos(x1_aw_deq_io_deq_bits_qos),
    .io_deq_bits_echo_tl_state_source(x1_aw_deq_io_deq_bits_echo_tl_state_source)
  );
  Queue_7 x1_w_deq ( // @[Decoupled.scala 375:21]
    .clock(x1_w_deq_clock),
    .reset(x1_w_deq_reset),
    .io_enq_ready(x1_w_deq_io_enq_ready),
    .io_enq_valid(x1_w_deq_io_enq_valid),
    .io_enq_bits_data(x1_w_deq_io_enq_bits_data),
    .io_enq_bits_strb(x1_w_deq_io_enq_bits_strb),
    .io_enq_bits_last(x1_w_deq_io_enq_bits_last),
    .io_deq_ready(x1_w_deq_io_deq_ready),
    .io_deq_valid(x1_w_deq_io_deq_valid),
    .io_deq_bits_data(x1_w_deq_io_deq_bits_data),
    .io_deq_bits_strb(x1_w_deq_io_deq_bits_strb),
    .io_deq_bits_last(x1_w_deq_io_deq_bits_last)
  );
  Queue_8 bundleIn_0_b_deq ( // @[Decoupled.scala 375:21]
    .clock(bundleIn_0_b_deq_clock),
    .reset(bundleIn_0_b_deq_reset),
    .io_enq_ready(bundleIn_0_b_deq_io_enq_ready),
    .io_enq_valid(bundleIn_0_b_deq_io_enq_valid),
    .io_enq_bits_id(bundleIn_0_b_deq_io_enq_bits_id),
    .io_enq_bits_echo_tl_state_source(bundleIn_0_b_deq_io_enq_bits_echo_tl_state_source),
    .io_deq_ready(bundleIn_0_b_deq_io_deq_ready),
    .io_deq_valid(bundleIn_0_b_deq_io_deq_valid),
    .io_deq_bits_id(bundleIn_0_b_deq_io_deq_bits_id),
    .io_deq_bits_echo_tl_state_source(bundleIn_0_b_deq_io_deq_bits_echo_tl_state_source)
  );
  Queue_6 x1_ar_deq ( // @[Decoupled.scala 375:21]
    .clock(x1_ar_deq_clock),
    .reset(x1_ar_deq_reset),
    .io_enq_ready(x1_ar_deq_io_enq_ready),
    .io_enq_valid(x1_ar_deq_io_enq_valid),
    .io_enq_bits_id(x1_ar_deq_io_enq_bits_id),
    .io_enq_bits_addr(x1_ar_deq_io_enq_bits_addr),
    .io_enq_bits_len(x1_ar_deq_io_enq_bits_len),
    .io_enq_bits_size(x1_ar_deq_io_enq_bits_size),
    .io_enq_bits_burst(x1_ar_deq_io_enq_bits_burst),
    .io_enq_bits_lock(x1_ar_deq_io_enq_bits_lock),
    .io_enq_bits_cache(x1_ar_deq_io_enq_bits_cache),
    .io_enq_bits_prot(x1_ar_deq_io_enq_bits_prot),
    .io_enq_bits_qos(x1_ar_deq_io_enq_bits_qos),
    .io_enq_bits_echo_tl_state_source(x1_ar_deq_io_enq_bits_echo_tl_state_source),
    .io_deq_ready(x1_ar_deq_io_deq_ready),
    .io_deq_valid(x1_ar_deq_io_deq_valid),
    .io_deq_bits_id(x1_ar_deq_io_deq_bits_id),
    .io_deq_bits_addr(x1_ar_deq_io_deq_bits_addr),
    .io_deq_bits_len(x1_ar_deq_io_deq_bits_len),
    .io_deq_bits_size(x1_ar_deq_io_deq_bits_size),
    .io_deq_bits_burst(x1_ar_deq_io_deq_bits_burst),
    .io_deq_bits_lock(x1_ar_deq_io_deq_bits_lock),
    .io_deq_bits_cache(x1_ar_deq_io_deq_bits_cache),
    .io_deq_bits_prot(x1_ar_deq_io_deq_bits_prot),
    .io_deq_bits_qos(x1_ar_deq_io_deq_bits_qos),
    .io_deq_bits_echo_tl_state_source(x1_ar_deq_io_deq_bits_echo_tl_state_source)
  );
  Queue_10 bundleIn_0_r_deq ( // @[Decoupled.scala 375:21]
    .clock(bundleIn_0_r_deq_clock),
    .reset(bundleIn_0_r_deq_reset),
    .io_enq_ready(bundleIn_0_r_deq_io_enq_ready),
    .io_enq_valid(bundleIn_0_r_deq_io_enq_valid),
    .io_enq_bits_id(bundleIn_0_r_deq_io_enq_bits_id),
    .io_enq_bits_data(bundleIn_0_r_deq_io_enq_bits_data),
    .io_enq_bits_echo_tl_state_source(bundleIn_0_r_deq_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(bundleIn_0_r_deq_io_enq_bits_last),
    .io_deq_ready(bundleIn_0_r_deq_io_deq_ready),
    .io_deq_valid(bundleIn_0_r_deq_io_deq_valid),
    .io_deq_bits_id(bundleIn_0_r_deq_io_deq_bits_id),
    .io_deq_bits_data(bundleIn_0_r_deq_io_deq_bits_data),
    .io_deq_bits_echo_tl_state_source(bundleIn_0_r_deq_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(bundleIn_0_r_deq_io_deq_bits_last)
  );
  assign auto_in_aw_ready = x1_aw_deq_io_enq_ready; // @[Nodes.scala 1215:84 Decoupled.scala 379:17]
  assign auto_in_w_ready = x1_w_deq_io_enq_ready; // @[Nodes.scala 1215:84 Decoupled.scala 379:17]
  assign auto_in_b_valid = bundleIn_0_b_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_in_b_bits_id = bundleIn_0_b_deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_b_bits_echo_tl_state_source = bundleIn_0_b_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_ar_ready = x1_ar_deq_io_enq_ready; // @[Nodes.scala 1215:84 Decoupled.scala 379:17]
  assign auto_in_r_valid = bundleIn_0_r_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_in_r_bits_id = bundleIn_0_r_deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_r_bits_data = bundleIn_0_r_deq_io_deq_bits_data; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_r_bits_echo_tl_state_source = bundleIn_0_r_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_r_bits_last = bundleIn_0_r_deq_io_deq_bits_last; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_valid = x1_aw_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_out_aw_bits_id = x1_aw_deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_addr = x1_aw_deq_io_deq_bits_addr; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_len = x1_aw_deq_io_deq_bits_len; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_size = x1_aw_deq_io_deq_bits_size; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_burst = x1_aw_deq_io_deq_bits_burst; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_lock = x1_aw_deq_io_deq_bits_lock; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_cache = x1_aw_deq_io_deq_bits_cache; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_prot = x1_aw_deq_io_deq_bits_prot; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_qos = x1_aw_deq_io_deq_bits_qos; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_echo_tl_state_source = x1_aw_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_w_valid = x1_w_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_out_w_bits_data = x1_w_deq_io_deq_bits_data; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_w_bits_strb = x1_w_deq_io_deq_bits_strb; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_w_bits_last = x1_w_deq_io_deq_bits_last; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_b_ready = bundleIn_0_b_deq_io_enq_ready; // @[Nodes.scala 1212:84 Decoupled.scala 379:17]
  assign auto_out_ar_valid = x1_ar_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_out_ar_bits_id = x1_ar_deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_addr = x1_ar_deq_io_deq_bits_addr; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_len = x1_ar_deq_io_deq_bits_len; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_size = x1_ar_deq_io_deq_bits_size; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_burst = x1_ar_deq_io_deq_bits_burst; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_lock = x1_ar_deq_io_deq_bits_lock; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_cache = x1_ar_deq_io_deq_bits_cache; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_prot = x1_ar_deq_io_deq_bits_prot; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_qos = x1_ar_deq_io_deq_bits_qos; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_echo_tl_state_source = x1_ar_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_r_ready = bundleIn_0_r_deq_io_enq_ready; // @[Nodes.scala 1212:84 Decoupled.scala 379:17]
  assign x1_aw_deq_clock = clock;
  assign x1_aw_deq_reset = reset;
  assign x1_aw_deq_io_enq_valid = auto_in_aw_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_id = auto_in_aw_bits_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_addr = auto_in_aw_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_len = auto_in_aw_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_size = auto_in_aw_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_burst = auto_in_aw_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_lock = auto_in_aw_bits_lock; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_cache = auto_in_aw_bits_cache; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_prot = auto_in_aw_bits_prot; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_qos = auto_in_aw_bits_qos; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_echo_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_deq_ready = auto_out_aw_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign x1_w_deq_clock = clock;
  assign x1_w_deq_reset = reset;
  assign x1_w_deq_io_enq_valid = auto_in_w_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_w_deq_io_enq_bits_data = auto_in_w_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_w_deq_io_enq_bits_strb = auto_in_w_bits_strb; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_w_deq_io_enq_bits_last = auto_in_w_bits_last; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_w_deq_io_deq_ready = auto_out_w_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_b_deq_clock = clock;
  assign bundleIn_0_b_deq_reset = reset;
  assign bundleIn_0_b_deq_io_enq_valid = auto_out_b_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_b_deq_io_enq_bits_id = auto_out_b_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_b_deq_io_enq_bits_echo_tl_state_source = auto_out_b_bits_echo_tl_state_source; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_b_deq_io_deq_ready = auto_in_b_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_clock = clock;
  assign x1_ar_deq_reset = reset;
  assign x1_ar_deq_io_enq_valid = auto_in_ar_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_id = auto_in_ar_bits_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_addr = auto_in_ar_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_len = auto_in_ar_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_size = auto_in_ar_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_burst = auto_in_ar_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_lock = auto_in_ar_bits_lock; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_cache = auto_in_ar_bits_cache; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_prot = auto_in_ar_bits_prot; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_qos = auto_in_ar_bits_qos; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_echo_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_deq_ready = auto_out_ar_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_clock = clock;
  assign bundleIn_0_r_deq_reset = reset;
  assign bundleIn_0_r_deq_io_enq_valid = auto_out_r_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_enq_bits_id = auto_out_r_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_enq_bits_data = auto_out_r_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_enq_bits_echo_tl_state_source = auto_out_r_bits_echo_tl_state_source; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_enq_bits_last = auto_out_r_bits_last; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_deq_ready = auto_in_r_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
endmodule
module Queue_16(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [511:0] io_enq_bits_data,
  input  [63:0]  io_enq_bits_strb,
  input          io_deq_ready,
  output         io_deq_valid,
  output [511:0] io_deq_bits_data,
  output [63:0]  io_deq_bits_strb,
  output         io_deq_bits_last
);
  reg [511:0] ram_data [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [511:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [511:0] ram_data_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 273:95]
  reg [63:0] ram_strb [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_strb_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_strb_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [63:0] ram_strb_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [63:0] ram_strb_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_strb_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_strb_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_strb_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_last [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_en; // @[Decoupled.scala 273:95]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 278:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_11 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 318:26 280:27 318:35]
  wire  do_enq = empty ? _GEN_11 : _do_enq_T; // @[Decoupled.scala 315:17 280:27]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 315:17 317:14 281:27]
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = 1'h0;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = empty ? _GEN_11 : _do_enq_T;
  assign ram_strb_io_deq_bits_MPORT_en = 1'h1;
  assign ram_strb_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_strb_io_deq_bits_MPORT_data = ram_strb[ram_strb_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_strb_MPORT_data = io_enq_bits_strb;
  assign ram_strb_MPORT_addr = 1'h0;
  assign ram_strb_MPORT_mask = 1'h1;
  assign ram_strb_MPORT_en = empty ? _GEN_11 : _do_enq_T;
  assign ram_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_last_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_last_io_deq_bits_MPORT_data = ram_last[ram_last_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_last_MPORT_data = 1'h1;
  assign ram_last_MPORT_addr = 1'h0;
  assign ram_last_MPORT_mask = 1'h1;
  assign ram_last_MPORT_en = empty ? _GEN_11 : _do_enq_T;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 302:16 314:{24,39}]
  assign io_deq_bits_data = empty ? io_enq_bits_data : ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_strb = empty ? io_enq_bits_strb : ram_strb_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_last = empty | ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  always @(posedge clock) begin
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_strb_MPORT_en & ram_strb_MPORT_mask) begin
      ram_strb[ram_strb_MPORT_addr] <= ram_strb_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_last_MPORT_en & ram_last_MPORT_mask) begin
      ram_last[ram_last_MPORT_addr] <= ram_last_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      if (empty) begin // @[Decoupled.scala 315:17]
        if (io_deq_ready) begin // @[Decoupled.scala 318:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 318:35]
        end else begin
          maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
        end
      end else begin
        maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
      end
    end
  end
endmodule
module Queue_17(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [6:0]  io_enq_bits_id,
  input  [33:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_len,
  input  [2:0]  io_enq_bits_size,
  input  [6:0]  io_enq_bits_echo_tl_state_source,
  input         io_enq_bits_wen,
  input         io_deq_ready,
  output        io_deq_valid,
  output [6:0]  io_deq_bits_id,
  output [33:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_len,
  output [2:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_burst,
  output        io_deq_bits_lock,
  output [3:0]  io_deq_bits_cache,
  output [2:0]  io_deq_bits_prot,
  output [3:0]  io_deq_bits_qos,
  output [6:0]  io_deq_bits_echo_tl_state_source,
  output        io_deq_bits_wen
);
  reg [6:0] ram_id [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [6:0] ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [6:0] ram_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [33:0] ram_addr [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_addr_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_addr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [33:0] ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [33:0] ram_addr_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_addr_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_addr_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_addr_MPORT_en; // @[Decoupled.scala 273:95]
  reg [7:0] ram_len [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_len_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_len_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [7:0] ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [7:0] ram_len_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_len_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_len_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_len_MPORT_en; // @[Decoupled.scala 273:95]
  reg [2:0] ram_size [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_size_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_burst [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_burst_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_burst_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_burst_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_burst_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_burst_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_burst_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_lock [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_lock_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_lock_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_lock_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_lock_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_lock_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_lock_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_lock_MPORT_en; // @[Decoupled.scala 273:95]
  reg [3:0] ram_cache [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_cache_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_cache_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [3:0] ram_cache_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [3:0] ram_cache_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_cache_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_cache_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_cache_MPORT_en; // @[Decoupled.scala 273:95]
  reg [2:0] ram_prot [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_prot_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_prot_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [2:0] ram_prot_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_prot_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_prot_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_prot_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_prot_MPORT_en; // @[Decoupled.scala 273:95]
  reg [3:0] ram_qos [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_qos_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_qos_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [3:0] ram_qos_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [3:0] ram_qos_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_qos_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_qos_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_qos_MPORT_en; // @[Decoupled.scala 273:95]
  reg [6:0] ram_echo_tl_state_source [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [6:0] ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [6:0] ram_echo_tl_state_source_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_wen [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_wen_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_wen_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_wen_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_wen_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_wen_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_wen_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_wen_MPORT_en; // @[Decoupled.scala 273:95]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 278:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_20 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 318:26 280:27 318:35]
  wire  do_enq = empty ? _GEN_20 : _do_enq_T; // @[Decoupled.scala 315:17 280:27]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 315:17 317:14 281:27]
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = 1'h0;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = empty ? _GEN_20 : _do_enq_T;
  assign ram_addr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_addr_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = 1'h0;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = empty ? _GEN_20 : _do_enq_T;
  assign ram_len_io_deq_bits_MPORT_en = 1'h1;
  assign ram_len_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_len_io_deq_bits_MPORT_data = ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_len_MPORT_data = io_enq_bits_len;
  assign ram_len_MPORT_addr = 1'h0;
  assign ram_len_MPORT_mask = 1'h1;
  assign ram_len_MPORT_en = empty ? _GEN_20 : _do_enq_T;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = 1'h0;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = empty ? _GEN_20 : _do_enq_T;
  assign ram_burst_io_deq_bits_MPORT_en = 1'h1;
  assign ram_burst_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_burst_io_deq_bits_MPORT_data = ram_burst[ram_burst_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_burst_MPORT_data = 2'h1;
  assign ram_burst_MPORT_addr = 1'h0;
  assign ram_burst_MPORT_mask = 1'h1;
  assign ram_burst_MPORT_en = empty ? _GEN_20 : _do_enq_T;
  assign ram_lock_io_deq_bits_MPORT_en = 1'h1;
  assign ram_lock_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_lock_io_deq_bits_MPORT_data = ram_lock[ram_lock_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_lock_MPORT_data = 1'h0;
  assign ram_lock_MPORT_addr = 1'h0;
  assign ram_lock_MPORT_mask = 1'h1;
  assign ram_lock_MPORT_en = empty ? _GEN_20 : _do_enq_T;
  assign ram_cache_io_deq_bits_MPORT_en = 1'h1;
  assign ram_cache_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_cache_io_deq_bits_MPORT_data = ram_cache[ram_cache_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_cache_MPORT_data = 4'h0;
  assign ram_cache_MPORT_addr = 1'h0;
  assign ram_cache_MPORT_mask = 1'h1;
  assign ram_cache_MPORT_en = empty ? _GEN_20 : _do_enq_T;
  assign ram_prot_io_deq_bits_MPORT_en = 1'h1;
  assign ram_prot_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_prot_io_deq_bits_MPORT_data = ram_prot[ram_prot_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_prot_MPORT_data = 3'h1;
  assign ram_prot_MPORT_addr = 1'h0;
  assign ram_prot_MPORT_mask = 1'h1;
  assign ram_prot_MPORT_en = empty ? _GEN_20 : _do_enq_T;
  assign ram_qos_io_deq_bits_MPORT_en = 1'h1;
  assign ram_qos_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_qos_io_deq_bits_MPORT_data = ram_qos[ram_qos_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_qos_MPORT_data = 4'h0;
  assign ram_qos_MPORT_addr = 1'h0;
  assign ram_qos_MPORT_mask = 1'h1;
  assign ram_qos_MPORT_en = empty ? _GEN_20 : _do_enq_T;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_data =
    ram_echo_tl_state_source[ram_echo_tl_state_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_echo_tl_state_source_MPORT_data = io_enq_bits_echo_tl_state_source;
  assign ram_echo_tl_state_source_MPORT_addr = 1'h0;
  assign ram_echo_tl_state_source_MPORT_mask = 1'h1;
  assign ram_echo_tl_state_source_MPORT_en = empty ? _GEN_20 : _do_enq_T;
  assign ram_wen_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wen_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wen_io_deq_bits_MPORT_data = ram_wen[ram_wen_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_wen_MPORT_data = io_enq_bits_wen;
  assign ram_wen_MPORT_addr = 1'h0;
  assign ram_wen_MPORT_mask = 1'h1;
  assign ram_wen_MPORT_en = empty ? _GEN_20 : _do_enq_T;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 302:16 314:{24,39}]
  assign io_deq_bits_id = empty ? io_enq_bits_id : ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_addr = empty ? io_enq_bits_addr : ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_len = empty ? io_enq_bits_len : ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_size = empty ? io_enq_bits_size : ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_burst = empty ? 2'h1 : ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_lock = empty ? 1'h0 : ram_lock_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_cache = empty ? 4'h0 : ram_cache_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_prot = empty ? 3'h1 : ram_prot_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_qos = empty ? 4'h0 : ram_qos_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_echo_tl_state_source = empty ? io_enq_bits_echo_tl_state_source :
    ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_wen = empty ? io_enq_bits_wen : ram_wen_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_len_MPORT_en & ram_len_MPORT_mask) begin
      ram_len[ram_len_MPORT_addr] <= ram_len_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_burst_MPORT_en & ram_burst_MPORT_mask) begin
      ram_burst[ram_burst_MPORT_addr] <= ram_burst_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_lock_MPORT_en & ram_lock_MPORT_mask) begin
      ram_lock[ram_lock_MPORT_addr] <= ram_lock_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_cache_MPORT_en & ram_cache_MPORT_mask) begin
      ram_cache[ram_cache_MPORT_addr] <= ram_cache_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_prot_MPORT_en & ram_prot_MPORT_mask) begin
      ram_prot[ram_prot_MPORT_addr] <= ram_prot_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_qos_MPORT_en & ram_qos_MPORT_mask) begin
      ram_qos[ram_qos_MPORT_addr] <= ram_qos_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_echo_tl_state_source_MPORT_en & ram_echo_tl_state_source_MPORT_mask) begin
      ram_echo_tl_state_source[ram_echo_tl_state_source_MPORT_addr] <= ram_echo_tl_state_source_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_wen_MPORT_en & ram_wen_MPORT_mask) begin
      ram_wen[ram_wen_MPORT_addr] <= ram_wen_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      if (empty) begin // @[Decoupled.scala 315:17]
        if (io_deq_ready) begin // @[Decoupled.scala 318:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 318:35]
        end else begin
          maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
        end
      end else begin
        maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
      end
    end
  end
endmodule
module TLToAXI4(
  input          clock,
  input          reset,
  output         auto_in_a_ready,
  input          auto_in_a_valid,
  input  [2:0]   auto_in_a_bits_opcode,
  input  [2:0]   auto_in_a_bits_size,
  input  [6:0]   auto_in_a_bits_source,
  input  [33:0]  auto_in_a_bits_address,
  input  [63:0]  auto_in_a_bits_mask,
  input  [511:0] auto_in_a_bits_data,
  input          auto_in_d_ready,
  output         auto_in_d_valid,
  output [6:0]   auto_in_d_bits_source,
  output [511:0] auto_in_d_bits_data,
  input          auto_out_aw_ready,
  output         auto_out_aw_valid,
  output [6:0]   auto_out_aw_bits_id,
  output [33:0]  auto_out_aw_bits_addr,
  output [7:0]   auto_out_aw_bits_len,
  output [2:0]   auto_out_aw_bits_size,
  output [1:0]   auto_out_aw_bits_burst,
  output         auto_out_aw_bits_lock,
  output [3:0]   auto_out_aw_bits_cache,
  output [2:0]   auto_out_aw_bits_prot,
  output [3:0]   auto_out_aw_bits_qos,
  output [6:0]   auto_out_aw_bits_echo_tl_state_source,
  input          auto_out_w_ready,
  output         auto_out_w_valid,
  output [511:0] auto_out_w_bits_data,
  output [63:0]  auto_out_w_bits_strb,
  output         auto_out_w_bits_last,
  output         auto_out_b_ready,
  input          auto_out_b_valid,
  input  [6:0]   auto_out_b_bits_id,
  input  [6:0]   auto_out_b_bits_echo_tl_state_source,
  input          auto_out_ar_ready,
  output         auto_out_ar_valid,
  output [6:0]   auto_out_ar_bits_id,
  output [33:0]  auto_out_ar_bits_addr,
  output [7:0]   auto_out_ar_bits_len,
  output [2:0]   auto_out_ar_bits_size,
  output [1:0]   auto_out_ar_bits_burst,
  output         auto_out_ar_bits_lock,
  output [3:0]   auto_out_ar_bits_cache,
  output [2:0]   auto_out_ar_bits_prot,
  output [3:0]   auto_out_ar_bits_qos,
  output [6:0]   auto_out_ar_bits_echo_tl_state_source,
  output         auto_out_r_ready,
  input          auto_out_r_valid,
  input  [6:0]   auto_out_r_bits_id,
  input  [511:0] auto_out_r_bits_data,
  input  [6:0]   auto_out_r_bits_echo_tl_state_source,
  input          auto_out_r_bits_last
);
  wire  deq_clock; // @[Decoupled.scala 375:21]
  wire  deq_reset; // @[Decoupled.scala 375:21]
  wire  deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [511:0] deq_io_enq_bits_data; // @[Decoupled.scala 375:21]
  wire [63:0] deq_io_enq_bits_strb; // @[Decoupled.scala 375:21]
  wire  deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [511:0] deq_io_deq_bits_data; // @[Decoupled.scala 375:21]
  wire [63:0] deq_io_deq_bits_strb; // @[Decoupled.scala 375:21]
  wire  deq_io_deq_bits_last; // @[Decoupled.scala 375:21]
  wire  queue_arw_deq_clock; // @[Decoupled.scala 375:21]
  wire  queue_arw_deq_reset; // @[Decoupled.scala 375:21]
  wire  queue_arw_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  queue_arw_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [6:0] queue_arw_deq_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire [33:0] queue_arw_deq_io_enq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] queue_arw_deq_io_enq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] queue_arw_deq_io_enq_bits_size; // @[Decoupled.scala 375:21]
  wire [6:0] queue_arw_deq_io_enq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire  queue_arw_deq_io_enq_bits_wen; // @[Decoupled.scala 375:21]
  wire  queue_arw_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  queue_arw_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [6:0] queue_arw_deq_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [33:0] queue_arw_deq_io_deq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] queue_arw_deq_io_deq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] queue_arw_deq_io_deq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] queue_arw_deq_io_deq_bits_burst; // @[Decoupled.scala 375:21]
  wire  queue_arw_deq_io_deq_bits_lock; // @[Decoupled.scala 375:21]
  wire [3:0] queue_arw_deq_io_deq_bits_cache; // @[Decoupled.scala 375:21]
  wire [2:0] queue_arw_deq_io_deq_bits_prot; // @[Decoupled.scala 375:21]
  wire [3:0] queue_arw_deq_io_deq_bits_qos; // @[Decoupled.scala 375:21]
  wire [6:0] queue_arw_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire  queue_arw_deq_io_deq_bits_wen; // @[Decoupled.scala 375:21]
  wire  a_isPut = ~auto_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  reg  count_66; // @[ToAXI4.scala 257:28]
  wire  idle_65 = ~count_66; // @[ToAXI4.scala 259:26]
  reg  count_65; // @[ToAXI4.scala 257:28]
  wire  idle_64 = ~count_65; // @[ToAXI4.scala 259:26]
  reg  count_64; // @[ToAXI4.scala 257:28]
  wire  idle_63 = ~count_64; // @[ToAXI4.scala 259:26]
  reg  count_63; // @[ToAXI4.scala 257:28]
  wire  idle_62 = ~count_63; // @[ToAXI4.scala 259:26]
  reg  count_62; // @[ToAXI4.scala 257:28]
  wire  idle_61 = ~count_62; // @[ToAXI4.scala 259:26]
  reg  count_61; // @[ToAXI4.scala 257:28]
  wire  idle_60 = ~count_61; // @[ToAXI4.scala 259:26]
  reg  count_60; // @[ToAXI4.scala 257:28]
  wire  idle_59 = ~count_60; // @[ToAXI4.scala 259:26]
  reg  count_59; // @[ToAXI4.scala 257:28]
  wire  idle_58 = ~count_59; // @[ToAXI4.scala 259:26]
  reg  count_58; // @[ToAXI4.scala 257:28]
  wire  idle_57 = ~count_58; // @[ToAXI4.scala 259:26]
  reg  count_57; // @[ToAXI4.scala 257:28]
  wire  idle_56 = ~count_57; // @[ToAXI4.scala 259:26]
  reg  count_56; // @[ToAXI4.scala 257:28]
  wire  idle_55 = ~count_56; // @[ToAXI4.scala 259:26]
  reg  count_55; // @[ToAXI4.scala 257:28]
  wire  idle_54 = ~count_55; // @[ToAXI4.scala 259:26]
  reg  count_54; // @[ToAXI4.scala 257:28]
  wire  idle_53 = ~count_54; // @[ToAXI4.scala 259:26]
  reg  count_53; // @[ToAXI4.scala 257:28]
  wire  idle_52 = ~count_53; // @[ToAXI4.scala 259:26]
  reg  count_52; // @[ToAXI4.scala 257:28]
  wire  idle_51 = ~count_52; // @[ToAXI4.scala 259:26]
  reg  count_51; // @[ToAXI4.scala 257:28]
  wire  idle_50 = ~count_51; // @[ToAXI4.scala 259:26]
  reg  count_50; // @[ToAXI4.scala 257:28]
  wire  idle_49 = ~count_50; // @[ToAXI4.scala 259:26]
  reg  count_49; // @[ToAXI4.scala 257:28]
  wire  idle_48 = ~count_49; // @[ToAXI4.scala 259:26]
  reg  count_48; // @[ToAXI4.scala 257:28]
  wire  idle_47 = ~count_48; // @[ToAXI4.scala 259:26]
  reg  count_47; // @[ToAXI4.scala 257:28]
  wire  idle_46 = ~count_47; // @[ToAXI4.scala 259:26]
  reg  count_46; // @[ToAXI4.scala 257:28]
  wire  idle_45 = ~count_46; // @[ToAXI4.scala 259:26]
  reg  count_45; // @[ToAXI4.scala 257:28]
  wire  idle_44 = ~count_45; // @[ToAXI4.scala 259:26]
  reg  count_44; // @[ToAXI4.scala 257:28]
  wire  idle_43 = ~count_44; // @[ToAXI4.scala 259:26]
  reg  count_43; // @[ToAXI4.scala 257:28]
  wire  idle_42 = ~count_43; // @[ToAXI4.scala 259:26]
  reg  count_42; // @[ToAXI4.scala 257:28]
  wire  idle_41 = ~count_42; // @[ToAXI4.scala 259:26]
  reg  count_41; // @[ToAXI4.scala 257:28]
  wire  idle_40 = ~count_41; // @[ToAXI4.scala 259:26]
  reg  count_40; // @[ToAXI4.scala 257:28]
  wire  idle_39 = ~count_40; // @[ToAXI4.scala 259:26]
  reg  count_39; // @[ToAXI4.scala 257:28]
  wire  idle_38 = ~count_39; // @[ToAXI4.scala 259:26]
  reg  count_38; // @[ToAXI4.scala 257:28]
  wire  idle_37 = ~count_38; // @[ToAXI4.scala 259:26]
  reg  count_37; // @[ToAXI4.scala 257:28]
  wire  idle_36 = ~count_37; // @[ToAXI4.scala 259:26]
  reg  count_36; // @[ToAXI4.scala 257:28]
  wire  idle_35 = ~count_36; // @[ToAXI4.scala 259:26]
  reg  count_35; // @[ToAXI4.scala 257:28]
  wire  idle_34 = ~count_35; // @[ToAXI4.scala 259:26]
  reg  count_34; // @[ToAXI4.scala 257:28]
  wire  idle_33 = ~count_34; // @[ToAXI4.scala 259:26]
  reg  count_33; // @[ToAXI4.scala 257:28]
  wire  idle_32 = ~count_33; // @[ToAXI4.scala 259:26]
  reg  count_32; // @[ToAXI4.scala 257:28]
  wire  idle_31 = ~count_32; // @[ToAXI4.scala 259:26]
  reg  count_31; // @[ToAXI4.scala 257:28]
  wire  idle_30 = ~count_31; // @[ToAXI4.scala 259:26]
  reg  count_30; // @[ToAXI4.scala 257:28]
  wire  idle_29 = ~count_30; // @[ToAXI4.scala 259:26]
  reg  count_29; // @[ToAXI4.scala 257:28]
  wire  idle_28 = ~count_29; // @[ToAXI4.scala 259:26]
  reg  count_28; // @[ToAXI4.scala 257:28]
  wire  idle_27 = ~count_28; // @[ToAXI4.scala 259:26]
  reg  count_27; // @[ToAXI4.scala 257:28]
  wire  idle_26 = ~count_27; // @[ToAXI4.scala 259:26]
  reg  count_26; // @[ToAXI4.scala 257:28]
  wire  idle_25 = ~count_26; // @[ToAXI4.scala 259:26]
  reg  count_25; // @[ToAXI4.scala 257:28]
  wire  idle_24 = ~count_25; // @[ToAXI4.scala 259:26]
  reg  count_24; // @[ToAXI4.scala 257:28]
  wire  idle_23 = ~count_24; // @[ToAXI4.scala 259:26]
  reg  count_23; // @[ToAXI4.scala 257:28]
  wire  idle_22 = ~count_23; // @[ToAXI4.scala 259:26]
  reg  count_22; // @[ToAXI4.scala 257:28]
  wire  idle_21 = ~count_22; // @[ToAXI4.scala 259:26]
  reg  count_21; // @[ToAXI4.scala 257:28]
  wire  idle_20 = ~count_21; // @[ToAXI4.scala 259:26]
  reg  count_20; // @[ToAXI4.scala 257:28]
  wire  idle_19 = ~count_20; // @[ToAXI4.scala 259:26]
  reg  count_19; // @[ToAXI4.scala 257:28]
  wire  idle_18 = ~count_19; // @[ToAXI4.scala 259:26]
  reg  count_18; // @[ToAXI4.scala 257:28]
  wire  idle_17 = ~count_18; // @[ToAXI4.scala 259:26]
  reg  count_17; // @[ToAXI4.scala 257:28]
  wire  idle_16 = ~count_17; // @[ToAXI4.scala 259:26]
  reg  count_16; // @[ToAXI4.scala 257:28]
  wire  idle_15 = ~count_16; // @[ToAXI4.scala 259:26]
  reg  count_15; // @[ToAXI4.scala 257:28]
  wire  idle_14 = ~count_15; // @[ToAXI4.scala 259:26]
  reg  count_14; // @[ToAXI4.scala 257:28]
  wire  idle_13 = ~count_14; // @[ToAXI4.scala 259:26]
  reg  count_13; // @[ToAXI4.scala 257:28]
  wire  idle_12 = ~count_13; // @[ToAXI4.scala 259:26]
  reg  count_12; // @[ToAXI4.scala 257:28]
  wire  idle_11 = ~count_12; // @[ToAXI4.scala 259:26]
  reg  count_11; // @[ToAXI4.scala 257:28]
  wire  idle_10 = ~count_11; // @[ToAXI4.scala 259:26]
  reg  count_10; // @[ToAXI4.scala 257:28]
  wire  idle_9 = ~count_10; // @[ToAXI4.scala 259:26]
  reg  count_9; // @[ToAXI4.scala 257:28]
  wire  idle_8 = ~count_9; // @[ToAXI4.scala 259:26]
  reg  count_8; // @[ToAXI4.scala 257:28]
  wire  idle_7 = ~count_8; // @[ToAXI4.scala 259:26]
  reg  count_7; // @[ToAXI4.scala 257:28]
  wire  idle_6 = ~count_7; // @[ToAXI4.scala 259:26]
  reg  count_6; // @[ToAXI4.scala 257:28]
  wire  idle_5 = ~count_6; // @[ToAXI4.scala 259:26]
  reg  count_5; // @[ToAXI4.scala 257:28]
  wire  idle_4 = ~count_5; // @[ToAXI4.scala 259:26]
  reg  count_4; // @[ToAXI4.scala 257:28]
  wire  idle_3 = ~count_4; // @[ToAXI4.scala 259:26]
  reg  count_3; // @[ToAXI4.scala 257:28]
  wire  idle_2 = ~count_3; // @[ToAXI4.scala 259:26]
  reg  count_2; // @[ToAXI4.scala 257:28]
  wire  idle_1 = ~count_2; // @[ToAXI4.scala 259:26]
  reg  count_1; // @[ToAXI4.scala 257:28]
  wire  idle = ~count_1; // @[ToAXI4.scala 259:26]
  wire  _GEN_69 = 7'h1 == auto_in_a_bits_source ? count_2 : count_1; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_70 = 7'h2 == auto_in_a_bits_source ? count_3 : _GEN_69; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_71 = 7'h3 == auto_in_a_bits_source ? count_4 : _GEN_70; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_72 = 7'h4 == auto_in_a_bits_source ? count_5 : _GEN_71; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_73 = 7'h5 == auto_in_a_bits_source ? count_6 : _GEN_72; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_74 = 7'h6 == auto_in_a_bits_source ? count_7 : _GEN_73; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_75 = 7'h7 == auto_in_a_bits_source ? count_8 : _GEN_74; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_76 = 7'h8 == auto_in_a_bits_source ? count_9 : _GEN_75; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_77 = 7'h9 == auto_in_a_bits_source ? count_10 : _GEN_76; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_78 = 7'ha == auto_in_a_bits_source ? count_11 : _GEN_77; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_79 = 7'hb == auto_in_a_bits_source ? count_12 : _GEN_78; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_80 = 7'hc == auto_in_a_bits_source ? count_13 : _GEN_79; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_81 = 7'hd == auto_in_a_bits_source ? count_14 : _GEN_80; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_82 = 7'he == auto_in_a_bits_source ? count_15 : _GEN_81; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_83 = 7'hf == auto_in_a_bits_source ? count_16 : _GEN_82; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_84 = 7'h10 == auto_in_a_bits_source ? count_17 : _GEN_83; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_85 = 7'h11 == auto_in_a_bits_source ? count_18 : _GEN_84; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_86 = 7'h12 == auto_in_a_bits_source ? count_19 : _GEN_85; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_87 = 7'h13 == auto_in_a_bits_source ? count_20 : _GEN_86; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_88 = 7'h14 == auto_in_a_bits_source ? count_21 : _GEN_87; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_89 = 7'h15 == auto_in_a_bits_source ? count_22 : _GEN_88; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_90 = 7'h16 == auto_in_a_bits_source ? count_23 : _GEN_89; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_91 = 7'h17 == auto_in_a_bits_source ? count_24 : _GEN_90; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_92 = 7'h18 == auto_in_a_bits_source ? count_25 : _GEN_91; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_93 = 7'h19 == auto_in_a_bits_source ? count_26 : _GEN_92; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_94 = 7'h1a == auto_in_a_bits_source ? count_27 : _GEN_93; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_95 = 7'h1b == auto_in_a_bits_source ? count_28 : _GEN_94; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_96 = 7'h1c == auto_in_a_bits_source ? count_29 : _GEN_95; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_97 = 7'h1d == auto_in_a_bits_source ? count_30 : _GEN_96; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_98 = 7'h1e == auto_in_a_bits_source ? count_31 : _GEN_97; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_99 = 7'h1f == auto_in_a_bits_source ? count_32 : _GEN_98; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_100 = 7'h20 == auto_in_a_bits_source ? count_33 : _GEN_99; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_101 = 7'h21 == auto_in_a_bits_source ? count_34 : _GEN_100; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_102 = 7'h22 == auto_in_a_bits_source ? count_35 : _GEN_101; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_103 = 7'h23 == auto_in_a_bits_source ? count_36 : _GEN_102; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_104 = 7'h24 == auto_in_a_bits_source ? count_37 : _GEN_103; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_105 = 7'h25 == auto_in_a_bits_source ? count_38 : _GEN_104; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_106 = 7'h26 == auto_in_a_bits_source ? count_39 : _GEN_105; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_107 = 7'h27 == auto_in_a_bits_source ? count_40 : _GEN_106; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_108 = 7'h28 == auto_in_a_bits_source ? count_41 : _GEN_107; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_109 = 7'h29 == auto_in_a_bits_source ? count_42 : _GEN_108; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_110 = 7'h2a == auto_in_a_bits_source ? count_43 : _GEN_109; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_111 = 7'h2b == auto_in_a_bits_source ? count_44 : _GEN_110; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_112 = 7'h2c == auto_in_a_bits_source ? count_45 : _GEN_111; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_113 = 7'h2d == auto_in_a_bits_source ? count_46 : _GEN_112; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_114 = 7'h2e == auto_in_a_bits_source ? count_47 : _GEN_113; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_115 = 7'h2f == auto_in_a_bits_source ? count_48 : _GEN_114; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_116 = 7'h30 == auto_in_a_bits_source ? count_49 : _GEN_115; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_117 = 7'h31 == auto_in_a_bits_source ? count_50 : _GEN_116; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_118 = 7'h32 == auto_in_a_bits_source ? count_51 : _GEN_117; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_119 = 7'h33 == auto_in_a_bits_source ? count_52 : _GEN_118; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_120 = 7'h34 == auto_in_a_bits_source ? count_53 : _GEN_119; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_121 = 7'h35 == auto_in_a_bits_source ? count_54 : _GEN_120; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_122 = 7'h36 == auto_in_a_bits_source ? count_55 : _GEN_121; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_123 = 7'h37 == auto_in_a_bits_source ? count_56 : _GEN_122; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_124 = 7'h38 == auto_in_a_bits_source ? count_57 : _GEN_123; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_125 = 7'h39 == auto_in_a_bits_source ? count_58 : _GEN_124; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_126 = 7'h3a == auto_in_a_bits_source ? count_59 : _GEN_125; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_127 = 7'h3b == auto_in_a_bits_source ? count_60 : _GEN_126; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_128 = 7'h3c == auto_in_a_bits_source ? count_61 : _GEN_127; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_129 = 7'h3d == auto_in_a_bits_source ? count_62 : _GEN_128; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_130 = 7'h3e == auto_in_a_bits_source ? count_63 : _GEN_129; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_131 = 7'h3f == auto_in_a_bits_source ? count_64 : _GEN_130; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_132 = 7'h40 == auto_in_a_bits_source ? count_65 : _GEN_131; // @[ToAXI4.scala 198:{49,49}]
  wire  _GEN_133 = 7'h41 == auto_in_a_bits_source ? count_66 : _GEN_132; // @[ToAXI4.scala 198:{49,49}]
  reg  counter; // @[Edges.scala 228:27]
  wire  a_first = ~counter; // @[Edges.scala 230:25]
  wire  stall = _GEN_133 & a_first; // @[ToAXI4.scala 198:49]
  wire  _bundleIn_0_a_ready_T = ~stall; // @[ToAXI4.scala 199:21]
  wire  out_arw_ready = queue_arw_deq_io_enq_ready; // @[ToAXI4.scala 150:25 Decoupled.scala 379:17]
  wire  out_w_ready = deq_io_enq_ready; // @[ToAXI4.scala 151:23 Decoupled.scala 379:17]
  wire  _bundleIn_0_a_ready_T_3 = a_isPut ? out_arw_ready & out_w_ready : out_arw_ready; // @[ToAXI4.scala 199:34]
  wire  bundleIn_0_a_ready = ~stall & _bundleIn_0_a_ready_T_3; // @[ToAXI4.scala 199:28]
  wire  done = bundleIn_0_a_ready & auto_in_a_valid; // @[Decoupled.scala 51:35]
  wire  counter1 = counter - 1'h1; // @[Edges.scala 229:28]
  wire  queue_arw_bits_wen = queue_arw_deq_io_deq_bits_wen; // @[Decoupled.scala 414:19 415:14]
  wire  queue_arw_valid = queue_arw_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  wire [6:0] _GEN_3 = 7'h1 == auto_in_a_bits_source ? 7'h1 : 7'h0; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_4 = 7'h2 == auto_in_a_bits_source ? 7'h2 : _GEN_3; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_5 = 7'h3 == auto_in_a_bits_source ? 7'h3 : _GEN_4; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_6 = 7'h4 == auto_in_a_bits_source ? 7'h4 : _GEN_5; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_7 = 7'h5 == auto_in_a_bits_source ? 7'h5 : _GEN_6; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_8 = 7'h6 == auto_in_a_bits_source ? 7'h6 : _GEN_7; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_9 = 7'h7 == auto_in_a_bits_source ? 7'h7 : _GEN_8; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_10 = 7'h8 == auto_in_a_bits_source ? 7'h8 : _GEN_9; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_11 = 7'h9 == auto_in_a_bits_source ? 7'h9 : _GEN_10; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_12 = 7'ha == auto_in_a_bits_source ? 7'ha : _GEN_11; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_13 = 7'hb == auto_in_a_bits_source ? 7'hb : _GEN_12; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_14 = 7'hc == auto_in_a_bits_source ? 7'hc : _GEN_13; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_15 = 7'hd == auto_in_a_bits_source ? 7'hd : _GEN_14; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_16 = 7'he == auto_in_a_bits_source ? 7'he : _GEN_15; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_17 = 7'hf == auto_in_a_bits_source ? 7'hf : _GEN_16; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_18 = 7'h10 == auto_in_a_bits_source ? 7'h10 : _GEN_17; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_19 = 7'h11 == auto_in_a_bits_source ? 7'h11 : _GEN_18; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_20 = 7'h12 == auto_in_a_bits_source ? 7'h12 : _GEN_19; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_21 = 7'h13 == auto_in_a_bits_source ? 7'h13 : _GEN_20; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_22 = 7'h14 == auto_in_a_bits_source ? 7'h14 : _GEN_21; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_23 = 7'h15 == auto_in_a_bits_source ? 7'h15 : _GEN_22; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_24 = 7'h16 == auto_in_a_bits_source ? 7'h16 : _GEN_23; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_25 = 7'h17 == auto_in_a_bits_source ? 7'h17 : _GEN_24; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_26 = 7'h18 == auto_in_a_bits_source ? 7'h18 : _GEN_25; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_27 = 7'h19 == auto_in_a_bits_source ? 7'h19 : _GEN_26; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_28 = 7'h1a == auto_in_a_bits_source ? 7'h1a : _GEN_27; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_29 = 7'h1b == auto_in_a_bits_source ? 7'h1b : _GEN_28; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_30 = 7'h1c == auto_in_a_bits_source ? 7'h1c : _GEN_29; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_31 = 7'h1d == auto_in_a_bits_source ? 7'h1d : _GEN_30; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_32 = 7'h1e == auto_in_a_bits_source ? 7'h1e : _GEN_31; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_33 = 7'h1f == auto_in_a_bits_source ? 7'h1f : _GEN_32; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_34 = 7'h20 == auto_in_a_bits_source ? 7'h20 : _GEN_33; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_35 = 7'h21 == auto_in_a_bits_source ? 7'h21 : _GEN_34; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_36 = 7'h22 == auto_in_a_bits_source ? 7'h22 : _GEN_35; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_37 = 7'h23 == auto_in_a_bits_source ? 7'h23 : _GEN_36; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_38 = 7'h24 == auto_in_a_bits_source ? 7'h24 : _GEN_37; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_39 = 7'h25 == auto_in_a_bits_source ? 7'h25 : _GEN_38; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_40 = 7'h26 == auto_in_a_bits_source ? 7'h26 : _GEN_39; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_41 = 7'h27 == auto_in_a_bits_source ? 7'h27 : _GEN_40; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_42 = 7'h28 == auto_in_a_bits_source ? 7'h28 : _GEN_41; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_43 = 7'h29 == auto_in_a_bits_source ? 7'h29 : _GEN_42; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_44 = 7'h2a == auto_in_a_bits_source ? 7'h2a : _GEN_43; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_45 = 7'h2b == auto_in_a_bits_source ? 7'h2b : _GEN_44; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_46 = 7'h2c == auto_in_a_bits_source ? 7'h2c : _GEN_45; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_47 = 7'h2d == auto_in_a_bits_source ? 7'h2d : _GEN_46; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_48 = 7'h2e == auto_in_a_bits_source ? 7'h2e : _GEN_47; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_49 = 7'h2f == auto_in_a_bits_source ? 7'h2f : _GEN_48; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_50 = 7'h30 == auto_in_a_bits_source ? 7'h30 : _GEN_49; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_51 = 7'h31 == auto_in_a_bits_source ? 7'h31 : _GEN_50; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_52 = 7'h32 == auto_in_a_bits_source ? 7'h32 : _GEN_51; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_53 = 7'h33 == auto_in_a_bits_source ? 7'h33 : _GEN_52; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_54 = 7'h34 == auto_in_a_bits_source ? 7'h34 : _GEN_53; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_55 = 7'h35 == auto_in_a_bits_source ? 7'h35 : _GEN_54; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_56 = 7'h36 == auto_in_a_bits_source ? 7'h36 : _GEN_55; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_57 = 7'h37 == auto_in_a_bits_source ? 7'h37 : _GEN_56; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_58 = 7'h38 == auto_in_a_bits_source ? 7'h38 : _GEN_57; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_59 = 7'h39 == auto_in_a_bits_source ? 7'h39 : _GEN_58; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_60 = 7'h3a == auto_in_a_bits_source ? 7'h3a : _GEN_59; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_61 = 7'h3b == auto_in_a_bits_source ? 7'h3b : _GEN_60; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_62 = 7'h3c == auto_in_a_bits_source ? 7'h3c : _GEN_61; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_63 = 7'h3d == auto_in_a_bits_source ? 7'h3d : _GEN_62; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_64 = 7'h3e == auto_in_a_bits_source ? 7'h3e : _GEN_63; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_65 = 7'h3f == auto_in_a_bits_source ? 7'h3f : _GEN_64; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] _GEN_66 = 7'h40 == auto_in_a_bits_source ? 7'h40 : _GEN_65; // @[ToAXI4.scala 169:{17,17}]
  wire [6:0] out_arw_bits_id = 7'h41 == auto_in_a_bits_source ? 7'h41 : _GEN_66; // @[ToAXI4.scala 169:{17,17}]
  wire [20:0] _out_arw_bits_len_T_1 = 21'h3fff << auto_in_a_bits_size; // @[package.scala 235:71]
  wire [13:0] _out_arw_bits_len_T_3 = ~_out_arw_bits_len_T_1[13:0]; // @[package.scala 235:46]
  wire  _out_arw_valid_T_1 = _bundleIn_0_a_ready_T & auto_in_a_valid; // @[ToAXI4.scala 200:31]
  wire  _out_arw_valid_T_4 = a_isPut ? out_w_ready : 1'h1; // @[ToAXI4.scala 200:51]
  wire  out_arw_valid = _bundleIn_0_a_ready_T & auto_in_a_valid & _out_arw_valid_T_4; // @[ToAXI4.scala 200:45]
  reg  r_holds_d; // @[ToAXI4.scala 209:30]
  reg [2:0] b_delay; // @[ToAXI4.scala 212:24]
  wire  r_wins = auto_out_r_valid & b_delay != 3'h7 | r_holds_d; // @[ToAXI4.scala 218:53]
  wire  x1_r_ready = auto_in_d_ready & r_wins; // @[ToAXI4.scala 220:33]
  wire  _T_2 = x1_r_ready & auto_out_r_valid; // @[Decoupled.scala 51:35]
  wire  x1_b_ready = auto_in_d_ready & ~r_wins; // @[ToAXI4.scala 221:33]
  wire [2:0] _b_delay_T_1 = b_delay + 3'h1; // @[ToAXI4.scala 214:28]
  wire  bundleIn_0_d_valid = r_wins ? auto_out_r_valid : auto_out_b_valid; // @[ToAXI4.scala 222:24]
  wire [127:0] _a_sel_T = 128'h1 << out_arw_bits_id; // @[OneHot.scala 64:12]
  wire  a_sel_0 = _a_sel_T[0]; // @[ToAXI4.scala 245:58]
  wire  a_sel_1 = _a_sel_T[1]; // @[ToAXI4.scala 245:58]
  wire  a_sel_2 = _a_sel_T[2]; // @[ToAXI4.scala 245:58]
  wire  a_sel_3 = _a_sel_T[3]; // @[ToAXI4.scala 245:58]
  wire  a_sel_4 = _a_sel_T[4]; // @[ToAXI4.scala 245:58]
  wire  a_sel_5 = _a_sel_T[5]; // @[ToAXI4.scala 245:58]
  wire  a_sel_6 = _a_sel_T[6]; // @[ToAXI4.scala 245:58]
  wire  a_sel_7 = _a_sel_T[7]; // @[ToAXI4.scala 245:58]
  wire  a_sel_8 = _a_sel_T[8]; // @[ToAXI4.scala 245:58]
  wire  a_sel_9 = _a_sel_T[9]; // @[ToAXI4.scala 245:58]
  wire  a_sel_10 = _a_sel_T[10]; // @[ToAXI4.scala 245:58]
  wire  a_sel_11 = _a_sel_T[11]; // @[ToAXI4.scala 245:58]
  wire  a_sel_12 = _a_sel_T[12]; // @[ToAXI4.scala 245:58]
  wire  a_sel_13 = _a_sel_T[13]; // @[ToAXI4.scala 245:58]
  wire  a_sel_14 = _a_sel_T[14]; // @[ToAXI4.scala 245:58]
  wire  a_sel_15 = _a_sel_T[15]; // @[ToAXI4.scala 245:58]
  wire  a_sel_16 = _a_sel_T[16]; // @[ToAXI4.scala 245:58]
  wire  a_sel_17 = _a_sel_T[17]; // @[ToAXI4.scala 245:58]
  wire  a_sel_18 = _a_sel_T[18]; // @[ToAXI4.scala 245:58]
  wire  a_sel_19 = _a_sel_T[19]; // @[ToAXI4.scala 245:58]
  wire  a_sel_20 = _a_sel_T[20]; // @[ToAXI4.scala 245:58]
  wire  a_sel_21 = _a_sel_T[21]; // @[ToAXI4.scala 245:58]
  wire  a_sel_22 = _a_sel_T[22]; // @[ToAXI4.scala 245:58]
  wire  a_sel_23 = _a_sel_T[23]; // @[ToAXI4.scala 245:58]
  wire  a_sel_24 = _a_sel_T[24]; // @[ToAXI4.scala 245:58]
  wire  a_sel_25 = _a_sel_T[25]; // @[ToAXI4.scala 245:58]
  wire  a_sel_26 = _a_sel_T[26]; // @[ToAXI4.scala 245:58]
  wire  a_sel_27 = _a_sel_T[27]; // @[ToAXI4.scala 245:58]
  wire  a_sel_28 = _a_sel_T[28]; // @[ToAXI4.scala 245:58]
  wire  a_sel_29 = _a_sel_T[29]; // @[ToAXI4.scala 245:58]
  wire  a_sel_30 = _a_sel_T[30]; // @[ToAXI4.scala 245:58]
  wire  a_sel_31 = _a_sel_T[31]; // @[ToAXI4.scala 245:58]
  wire  a_sel_32 = _a_sel_T[32]; // @[ToAXI4.scala 245:58]
  wire  a_sel_33 = _a_sel_T[33]; // @[ToAXI4.scala 245:58]
  wire  a_sel_34 = _a_sel_T[34]; // @[ToAXI4.scala 245:58]
  wire  a_sel_35 = _a_sel_T[35]; // @[ToAXI4.scala 245:58]
  wire  a_sel_36 = _a_sel_T[36]; // @[ToAXI4.scala 245:58]
  wire  a_sel_37 = _a_sel_T[37]; // @[ToAXI4.scala 245:58]
  wire  a_sel_38 = _a_sel_T[38]; // @[ToAXI4.scala 245:58]
  wire  a_sel_39 = _a_sel_T[39]; // @[ToAXI4.scala 245:58]
  wire  a_sel_40 = _a_sel_T[40]; // @[ToAXI4.scala 245:58]
  wire  a_sel_41 = _a_sel_T[41]; // @[ToAXI4.scala 245:58]
  wire  a_sel_42 = _a_sel_T[42]; // @[ToAXI4.scala 245:58]
  wire  a_sel_43 = _a_sel_T[43]; // @[ToAXI4.scala 245:58]
  wire  a_sel_44 = _a_sel_T[44]; // @[ToAXI4.scala 245:58]
  wire  a_sel_45 = _a_sel_T[45]; // @[ToAXI4.scala 245:58]
  wire  a_sel_46 = _a_sel_T[46]; // @[ToAXI4.scala 245:58]
  wire  a_sel_47 = _a_sel_T[47]; // @[ToAXI4.scala 245:58]
  wire  a_sel_48 = _a_sel_T[48]; // @[ToAXI4.scala 245:58]
  wire  a_sel_49 = _a_sel_T[49]; // @[ToAXI4.scala 245:58]
  wire  a_sel_50 = _a_sel_T[50]; // @[ToAXI4.scala 245:58]
  wire  a_sel_51 = _a_sel_T[51]; // @[ToAXI4.scala 245:58]
  wire  a_sel_52 = _a_sel_T[52]; // @[ToAXI4.scala 245:58]
  wire  a_sel_53 = _a_sel_T[53]; // @[ToAXI4.scala 245:58]
  wire  a_sel_54 = _a_sel_T[54]; // @[ToAXI4.scala 245:58]
  wire  a_sel_55 = _a_sel_T[55]; // @[ToAXI4.scala 245:58]
  wire  a_sel_56 = _a_sel_T[56]; // @[ToAXI4.scala 245:58]
  wire  a_sel_57 = _a_sel_T[57]; // @[ToAXI4.scala 245:58]
  wire  a_sel_58 = _a_sel_T[58]; // @[ToAXI4.scala 245:58]
  wire  a_sel_59 = _a_sel_T[59]; // @[ToAXI4.scala 245:58]
  wire  a_sel_60 = _a_sel_T[60]; // @[ToAXI4.scala 245:58]
  wire  a_sel_61 = _a_sel_T[61]; // @[ToAXI4.scala 245:58]
  wire  a_sel_62 = _a_sel_T[62]; // @[ToAXI4.scala 245:58]
  wire  a_sel_63 = _a_sel_T[63]; // @[ToAXI4.scala 245:58]
  wire  a_sel_64 = _a_sel_T[64]; // @[ToAXI4.scala 245:58]
  wire  a_sel_65 = _a_sel_T[65]; // @[ToAXI4.scala 245:58]
  wire [6:0] d_sel_shiftAmount = r_wins ? auto_out_r_bits_id : auto_out_b_bits_id; // @[ToAXI4.scala 246:31]
  wire [127:0] _d_sel_T_1 = 128'h1 << d_sel_shiftAmount; // @[OneHot.scala 64:12]
  wire  d_sel_0 = _d_sel_T_1[0]; // @[ToAXI4.scala 246:93]
  wire  d_sel_1 = _d_sel_T_1[1]; // @[ToAXI4.scala 246:93]
  wire  d_sel_2 = _d_sel_T_1[2]; // @[ToAXI4.scala 246:93]
  wire  d_sel_3 = _d_sel_T_1[3]; // @[ToAXI4.scala 246:93]
  wire  d_sel_4 = _d_sel_T_1[4]; // @[ToAXI4.scala 246:93]
  wire  d_sel_5 = _d_sel_T_1[5]; // @[ToAXI4.scala 246:93]
  wire  d_sel_6 = _d_sel_T_1[6]; // @[ToAXI4.scala 246:93]
  wire  d_sel_7 = _d_sel_T_1[7]; // @[ToAXI4.scala 246:93]
  wire  d_sel_8 = _d_sel_T_1[8]; // @[ToAXI4.scala 246:93]
  wire  d_sel_9 = _d_sel_T_1[9]; // @[ToAXI4.scala 246:93]
  wire  d_sel_10 = _d_sel_T_1[10]; // @[ToAXI4.scala 246:93]
  wire  d_sel_11 = _d_sel_T_1[11]; // @[ToAXI4.scala 246:93]
  wire  d_sel_12 = _d_sel_T_1[12]; // @[ToAXI4.scala 246:93]
  wire  d_sel_13 = _d_sel_T_1[13]; // @[ToAXI4.scala 246:93]
  wire  d_sel_14 = _d_sel_T_1[14]; // @[ToAXI4.scala 246:93]
  wire  d_sel_15 = _d_sel_T_1[15]; // @[ToAXI4.scala 246:93]
  wire  d_sel_16 = _d_sel_T_1[16]; // @[ToAXI4.scala 246:93]
  wire  d_sel_17 = _d_sel_T_1[17]; // @[ToAXI4.scala 246:93]
  wire  d_sel_18 = _d_sel_T_1[18]; // @[ToAXI4.scala 246:93]
  wire  d_sel_19 = _d_sel_T_1[19]; // @[ToAXI4.scala 246:93]
  wire  d_sel_20 = _d_sel_T_1[20]; // @[ToAXI4.scala 246:93]
  wire  d_sel_21 = _d_sel_T_1[21]; // @[ToAXI4.scala 246:93]
  wire  d_sel_22 = _d_sel_T_1[22]; // @[ToAXI4.scala 246:93]
  wire  d_sel_23 = _d_sel_T_1[23]; // @[ToAXI4.scala 246:93]
  wire  d_sel_24 = _d_sel_T_1[24]; // @[ToAXI4.scala 246:93]
  wire  d_sel_25 = _d_sel_T_1[25]; // @[ToAXI4.scala 246:93]
  wire  d_sel_26 = _d_sel_T_1[26]; // @[ToAXI4.scala 246:93]
  wire  d_sel_27 = _d_sel_T_1[27]; // @[ToAXI4.scala 246:93]
  wire  d_sel_28 = _d_sel_T_1[28]; // @[ToAXI4.scala 246:93]
  wire  d_sel_29 = _d_sel_T_1[29]; // @[ToAXI4.scala 246:93]
  wire  d_sel_30 = _d_sel_T_1[30]; // @[ToAXI4.scala 246:93]
  wire  d_sel_31 = _d_sel_T_1[31]; // @[ToAXI4.scala 246:93]
  wire  d_sel_32 = _d_sel_T_1[32]; // @[ToAXI4.scala 246:93]
  wire  d_sel_33 = _d_sel_T_1[33]; // @[ToAXI4.scala 246:93]
  wire  d_sel_34 = _d_sel_T_1[34]; // @[ToAXI4.scala 246:93]
  wire  d_sel_35 = _d_sel_T_1[35]; // @[ToAXI4.scala 246:93]
  wire  d_sel_36 = _d_sel_T_1[36]; // @[ToAXI4.scala 246:93]
  wire  d_sel_37 = _d_sel_T_1[37]; // @[ToAXI4.scala 246:93]
  wire  d_sel_38 = _d_sel_T_1[38]; // @[ToAXI4.scala 246:93]
  wire  d_sel_39 = _d_sel_T_1[39]; // @[ToAXI4.scala 246:93]
  wire  d_sel_40 = _d_sel_T_1[40]; // @[ToAXI4.scala 246:93]
  wire  d_sel_41 = _d_sel_T_1[41]; // @[ToAXI4.scala 246:93]
  wire  d_sel_42 = _d_sel_T_1[42]; // @[ToAXI4.scala 246:93]
  wire  d_sel_43 = _d_sel_T_1[43]; // @[ToAXI4.scala 246:93]
  wire  d_sel_44 = _d_sel_T_1[44]; // @[ToAXI4.scala 246:93]
  wire  d_sel_45 = _d_sel_T_1[45]; // @[ToAXI4.scala 246:93]
  wire  d_sel_46 = _d_sel_T_1[46]; // @[ToAXI4.scala 246:93]
  wire  d_sel_47 = _d_sel_T_1[47]; // @[ToAXI4.scala 246:93]
  wire  d_sel_48 = _d_sel_T_1[48]; // @[ToAXI4.scala 246:93]
  wire  d_sel_49 = _d_sel_T_1[49]; // @[ToAXI4.scala 246:93]
  wire  d_sel_50 = _d_sel_T_1[50]; // @[ToAXI4.scala 246:93]
  wire  d_sel_51 = _d_sel_T_1[51]; // @[ToAXI4.scala 246:93]
  wire  d_sel_52 = _d_sel_T_1[52]; // @[ToAXI4.scala 246:93]
  wire  d_sel_53 = _d_sel_T_1[53]; // @[ToAXI4.scala 246:93]
  wire  d_sel_54 = _d_sel_T_1[54]; // @[ToAXI4.scala 246:93]
  wire  d_sel_55 = _d_sel_T_1[55]; // @[ToAXI4.scala 246:93]
  wire  d_sel_56 = _d_sel_T_1[56]; // @[ToAXI4.scala 246:93]
  wire  d_sel_57 = _d_sel_T_1[57]; // @[ToAXI4.scala 246:93]
  wire  d_sel_58 = _d_sel_T_1[58]; // @[ToAXI4.scala 246:93]
  wire  d_sel_59 = _d_sel_T_1[59]; // @[ToAXI4.scala 246:93]
  wire  d_sel_60 = _d_sel_T_1[60]; // @[ToAXI4.scala 246:93]
  wire  d_sel_61 = _d_sel_T_1[61]; // @[ToAXI4.scala 246:93]
  wire  d_sel_62 = _d_sel_T_1[62]; // @[ToAXI4.scala 246:93]
  wire  d_sel_63 = _d_sel_T_1[63]; // @[ToAXI4.scala 246:93]
  wire  d_sel_64 = _d_sel_T_1[64]; // @[ToAXI4.scala 246:93]
  wire  d_sel_65 = _d_sel_T_1[65]; // @[ToAXI4.scala 246:93]
  wire  d_last = r_wins ? auto_out_r_bits_last : 1'h1; // @[ToAXI4.scala 247:23]
  wire  _inc_T = out_arw_ready & out_arw_valid; // @[Decoupled.scala 51:35]
  wire  inc = a_sel_0 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  _dec_T_1 = auto_in_d_ready & bundleIn_0_d_valid; // @[Decoupled.scala 51:35]
  wire  dec = d_sel_0 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_2 = count_1 + inc; // @[ToAXI4.scala 263:24]
  wire  _T_10 = ~reset; // @[ToAXI4.scala 265:16]
  wire  inc_1 = a_sel_1 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_1 = d_sel_1 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_6 = count_2 + inc_1; // @[ToAXI4.scala 263:24]
  wire  inc_2 = a_sel_2 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_2 = d_sel_2 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_10 = count_3 + inc_2; // @[ToAXI4.scala 263:24]
  wire  inc_3 = a_sel_3 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_3 = d_sel_3 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_14 = count_4 + inc_3; // @[ToAXI4.scala 263:24]
  wire  inc_4 = a_sel_4 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_4 = d_sel_4 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_18 = count_5 + inc_4; // @[ToAXI4.scala 263:24]
  wire  inc_5 = a_sel_5 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_5 = d_sel_5 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_22 = count_6 + inc_5; // @[ToAXI4.scala 263:24]
  wire  inc_6 = a_sel_6 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_6 = d_sel_6 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_26 = count_7 + inc_6; // @[ToAXI4.scala 263:24]
  wire  inc_7 = a_sel_7 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_7 = d_sel_7 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_30 = count_8 + inc_7; // @[ToAXI4.scala 263:24]
  wire  inc_8 = a_sel_8 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_8 = d_sel_8 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_34 = count_9 + inc_8; // @[ToAXI4.scala 263:24]
  wire  inc_9 = a_sel_9 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_9 = d_sel_9 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_38 = count_10 + inc_9; // @[ToAXI4.scala 263:24]
  wire  inc_10 = a_sel_10 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_10 = d_sel_10 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_42 = count_11 + inc_10; // @[ToAXI4.scala 263:24]
  wire  inc_11 = a_sel_11 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_11 = d_sel_11 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_46 = count_12 + inc_11; // @[ToAXI4.scala 263:24]
  wire  inc_12 = a_sel_12 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_12 = d_sel_12 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_50 = count_13 + inc_12; // @[ToAXI4.scala 263:24]
  wire  inc_13 = a_sel_13 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_13 = d_sel_13 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_54 = count_14 + inc_13; // @[ToAXI4.scala 263:24]
  wire  inc_14 = a_sel_14 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_14 = d_sel_14 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_58 = count_15 + inc_14; // @[ToAXI4.scala 263:24]
  wire  inc_15 = a_sel_15 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_15 = d_sel_15 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_62 = count_16 + inc_15; // @[ToAXI4.scala 263:24]
  wire  inc_16 = a_sel_16 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_16 = d_sel_16 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_66 = count_17 + inc_16; // @[ToAXI4.scala 263:24]
  wire  inc_17 = a_sel_17 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_17 = d_sel_17 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_70 = count_18 + inc_17; // @[ToAXI4.scala 263:24]
  wire  inc_18 = a_sel_18 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_18 = d_sel_18 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_74 = count_19 + inc_18; // @[ToAXI4.scala 263:24]
  wire  inc_19 = a_sel_19 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_19 = d_sel_19 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_78 = count_20 + inc_19; // @[ToAXI4.scala 263:24]
  wire  inc_20 = a_sel_20 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_20 = d_sel_20 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_82 = count_21 + inc_20; // @[ToAXI4.scala 263:24]
  wire  inc_21 = a_sel_21 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_21 = d_sel_21 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_86 = count_22 + inc_21; // @[ToAXI4.scala 263:24]
  wire  inc_22 = a_sel_22 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_22 = d_sel_22 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_90 = count_23 + inc_22; // @[ToAXI4.scala 263:24]
  wire  inc_23 = a_sel_23 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_23 = d_sel_23 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_94 = count_24 + inc_23; // @[ToAXI4.scala 263:24]
  wire  inc_24 = a_sel_24 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_24 = d_sel_24 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_98 = count_25 + inc_24; // @[ToAXI4.scala 263:24]
  wire  inc_25 = a_sel_25 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_25 = d_sel_25 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_102 = count_26 + inc_25; // @[ToAXI4.scala 263:24]
  wire  inc_26 = a_sel_26 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_26 = d_sel_26 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_106 = count_27 + inc_26; // @[ToAXI4.scala 263:24]
  wire  inc_27 = a_sel_27 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_27 = d_sel_27 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_110 = count_28 + inc_27; // @[ToAXI4.scala 263:24]
  wire  inc_28 = a_sel_28 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_28 = d_sel_28 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_114 = count_29 + inc_28; // @[ToAXI4.scala 263:24]
  wire  inc_29 = a_sel_29 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_29 = d_sel_29 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_118 = count_30 + inc_29; // @[ToAXI4.scala 263:24]
  wire  inc_30 = a_sel_30 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_30 = d_sel_30 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_122 = count_31 + inc_30; // @[ToAXI4.scala 263:24]
  wire  inc_31 = a_sel_31 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_31 = d_sel_31 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_126 = count_32 + inc_31; // @[ToAXI4.scala 263:24]
  wire  inc_32 = a_sel_32 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_32 = d_sel_32 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_130 = count_33 + inc_32; // @[ToAXI4.scala 263:24]
  wire  inc_33 = a_sel_33 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_33 = d_sel_33 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_134 = count_34 + inc_33; // @[ToAXI4.scala 263:24]
  wire  inc_34 = a_sel_34 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_34 = d_sel_34 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_138 = count_35 + inc_34; // @[ToAXI4.scala 263:24]
  wire  inc_35 = a_sel_35 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_35 = d_sel_35 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_142 = count_36 + inc_35; // @[ToAXI4.scala 263:24]
  wire  inc_36 = a_sel_36 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_36 = d_sel_36 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_146 = count_37 + inc_36; // @[ToAXI4.scala 263:24]
  wire  inc_37 = a_sel_37 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_37 = d_sel_37 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_150 = count_38 + inc_37; // @[ToAXI4.scala 263:24]
  wire  inc_38 = a_sel_38 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_38 = d_sel_38 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_154 = count_39 + inc_38; // @[ToAXI4.scala 263:24]
  wire  inc_39 = a_sel_39 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_39 = d_sel_39 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_158 = count_40 + inc_39; // @[ToAXI4.scala 263:24]
  wire  inc_40 = a_sel_40 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_40 = d_sel_40 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_162 = count_41 + inc_40; // @[ToAXI4.scala 263:24]
  wire  inc_41 = a_sel_41 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_41 = d_sel_41 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_166 = count_42 + inc_41; // @[ToAXI4.scala 263:24]
  wire  inc_42 = a_sel_42 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_42 = d_sel_42 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_170 = count_43 + inc_42; // @[ToAXI4.scala 263:24]
  wire  inc_43 = a_sel_43 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_43 = d_sel_43 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_174 = count_44 + inc_43; // @[ToAXI4.scala 263:24]
  wire  inc_44 = a_sel_44 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_44 = d_sel_44 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_178 = count_45 + inc_44; // @[ToAXI4.scala 263:24]
  wire  inc_45 = a_sel_45 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_45 = d_sel_45 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_182 = count_46 + inc_45; // @[ToAXI4.scala 263:24]
  wire  inc_46 = a_sel_46 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_46 = d_sel_46 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_186 = count_47 + inc_46; // @[ToAXI4.scala 263:24]
  wire  inc_47 = a_sel_47 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_47 = d_sel_47 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_190 = count_48 + inc_47; // @[ToAXI4.scala 263:24]
  wire  inc_48 = a_sel_48 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_48 = d_sel_48 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_194 = count_49 + inc_48; // @[ToAXI4.scala 263:24]
  wire  inc_49 = a_sel_49 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_49 = d_sel_49 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_198 = count_50 + inc_49; // @[ToAXI4.scala 263:24]
  wire  inc_50 = a_sel_50 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_50 = d_sel_50 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_202 = count_51 + inc_50; // @[ToAXI4.scala 263:24]
  wire  inc_51 = a_sel_51 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_51 = d_sel_51 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_206 = count_52 + inc_51; // @[ToAXI4.scala 263:24]
  wire  inc_52 = a_sel_52 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_52 = d_sel_52 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_210 = count_53 + inc_52; // @[ToAXI4.scala 263:24]
  wire  inc_53 = a_sel_53 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_53 = d_sel_53 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_214 = count_54 + inc_53; // @[ToAXI4.scala 263:24]
  wire  inc_54 = a_sel_54 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_54 = d_sel_54 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_218 = count_55 + inc_54; // @[ToAXI4.scala 263:24]
  wire  inc_55 = a_sel_55 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_55 = d_sel_55 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_222 = count_56 + inc_55; // @[ToAXI4.scala 263:24]
  wire  inc_56 = a_sel_56 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_56 = d_sel_56 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_226 = count_57 + inc_56; // @[ToAXI4.scala 263:24]
  wire  inc_57 = a_sel_57 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_57 = d_sel_57 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_230 = count_58 + inc_57; // @[ToAXI4.scala 263:24]
  wire  inc_58 = a_sel_58 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_58 = d_sel_58 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_234 = count_59 + inc_58; // @[ToAXI4.scala 263:24]
  wire  inc_59 = a_sel_59 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_59 = d_sel_59 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_238 = count_60 + inc_59; // @[ToAXI4.scala 263:24]
  wire  inc_60 = a_sel_60 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_60 = d_sel_60 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_242 = count_61 + inc_60; // @[ToAXI4.scala 263:24]
  wire  inc_61 = a_sel_61 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_61 = d_sel_61 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_246 = count_62 + inc_61; // @[ToAXI4.scala 263:24]
  wire  inc_62 = a_sel_62 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_62 = d_sel_62 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_250 = count_63 + inc_62; // @[ToAXI4.scala 263:24]
  wire  inc_63 = a_sel_63 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_63 = d_sel_63 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_254 = count_64 + inc_63; // @[ToAXI4.scala 263:24]
  wire  inc_64 = a_sel_64 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_64 = d_sel_64 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_258 = count_65 + inc_64; // @[ToAXI4.scala 263:24]
  wire  inc_65 = a_sel_65 & _inc_T; // @[ToAXI4.scala 261:22]
  wire  dec_65 = d_sel_65 & d_last & _dec_T_1; // @[ToAXI4.scala 262:32]
  wire  _count_T_262 = count_66 + inc_65; // @[ToAXI4.scala 263:24]
  Queue_16 deq ( // @[Decoupled.scala 375:21]
    .clock(deq_clock),
    .reset(deq_reset),
    .io_enq_ready(deq_io_enq_ready),
    .io_enq_valid(deq_io_enq_valid),
    .io_enq_bits_data(deq_io_enq_bits_data),
    .io_enq_bits_strb(deq_io_enq_bits_strb),
    .io_deq_ready(deq_io_deq_ready),
    .io_deq_valid(deq_io_deq_valid),
    .io_deq_bits_data(deq_io_deq_bits_data),
    .io_deq_bits_strb(deq_io_deq_bits_strb),
    .io_deq_bits_last(deq_io_deq_bits_last)
  );
  Queue_17 queue_arw_deq ( // @[Decoupled.scala 375:21]
    .clock(queue_arw_deq_clock),
    .reset(queue_arw_deq_reset),
    .io_enq_ready(queue_arw_deq_io_enq_ready),
    .io_enq_valid(queue_arw_deq_io_enq_valid),
    .io_enq_bits_id(queue_arw_deq_io_enq_bits_id),
    .io_enq_bits_addr(queue_arw_deq_io_enq_bits_addr),
    .io_enq_bits_len(queue_arw_deq_io_enq_bits_len),
    .io_enq_bits_size(queue_arw_deq_io_enq_bits_size),
    .io_enq_bits_echo_tl_state_source(queue_arw_deq_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_wen(queue_arw_deq_io_enq_bits_wen),
    .io_deq_ready(queue_arw_deq_io_deq_ready),
    .io_deq_valid(queue_arw_deq_io_deq_valid),
    .io_deq_bits_id(queue_arw_deq_io_deq_bits_id),
    .io_deq_bits_addr(queue_arw_deq_io_deq_bits_addr),
    .io_deq_bits_len(queue_arw_deq_io_deq_bits_len),
    .io_deq_bits_size(queue_arw_deq_io_deq_bits_size),
    .io_deq_bits_burst(queue_arw_deq_io_deq_bits_burst),
    .io_deq_bits_lock(queue_arw_deq_io_deq_bits_lock),
    .io_deq_bits_cache(queue_arw_deq_io_deq_bits_cache),
    .io_deq_bits_prot(queue_arw_deq_io_deq_bits_prot),
    .io_deq_bits_qos(queue_arw_deq_io_deq_bits_qos),
    .io_deq_bits_echo_tl_state_source(queue_arw_deq_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_wen(queue_arw_deq_io_deq_bits_wen)
  );
  assign auto_in_a_ready = ~stall & _bundleIn_0_a_ready_T_3; // @[ToAXI4.scala 199:28]
  assign auto_in_d_valid = r_wins ? auto_out_r_valid : auto_out_b_valid; // @[ToAXI4.scala 222:24]
  assign auto_in_d_bits_source = r_wins ? auto_out_r_bits_echo_tl_state_source : auto_out_b_bits_echo_tl_state_source; // @[ToAXI4.scala 240:23]
  assign auto_in_d_bits_data = auto_out_r_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_out_aw_valid = queue_arw_valid & queue_arw_bits_wen; // @[ToAXI4.scala 159:39]
  assign auto_out_aw_bits_id = queue_arw_deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_addr = queue_arw_deq_io_deq_bits_addr; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_len = queue_arw_deq_io_deq_bits_len; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_size = queue_arw_deq_io_deq_bits_size; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_burst = queue_arw_deq_io_deq_bits_burst; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_lock = queue_arw_deq_io_deq_bits_lock; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_cache = queue_arw_deq_io_deq_bits_cache; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_prot = queue_arw_deq_io_deq_bits_prot; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_qos = queue_arw_deq_io_deq_bits_qos; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_echo_tl_state_source = queue_arw_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_w_valid = deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_out_w_bits_data = deq_io_deq_bits_data; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_w_bits_strb = deq_io_deq_bits_strb; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_w_bits_last = deq_io_deq_bits_last; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_b_ready = auto_in_d_ready & ~r_wins; // @[ToAXI4.scala 221:33]
  assign auto_out_ar_valid = queue_arw_valid & ~queue_arw_bits_wen; // @[ToAXI4.scala 158:39]
  assign auto_out_ar_bits_id = queue_arw_deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_addr = queue_arw_deq_io_deq_bits_addr; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_len = queue_arw_deq_io_deq_bits_len; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_size = queue_arw_deq_io_deq_bits_size; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_burst = queue_arw_deq_io_deq_bits_burst; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_lock = queue_arw_deq_io_deq_bits_lock; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_cache = queue_arw_deq_io_deq_bits_cache; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_prot = queue_arw_deq_io_deq_bits_prot; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_qos = queue_arw_deq_io_deq_bits_qos; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_echo_tl_state_source = queue_arw_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_r_ready = auto_in_d_ready & r_wins; // @[ToAXI4.scala 220:33]
  assign deq_clock = clock;
  assign deq_reset = reset;
  assign deq_io_enq_valid = _out_arw_valid_T_1 & a_isPut & out_arw_ready; // @[ToAXI4.scala 202:54]
  assign deq_io_enq_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign deq_io_enq_bits_strb = auto_in_a_bits_mask; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign deq_io_deq_ready = auto_out_w_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign queue_arw_deq_clock = clock;
  assign queue_arw_deq_reset = reset;
  assign queue_arw_deq_io_enq_valid = _bundleIn_0_a_ready_T & auto_in_a_valid & _out_arw_valid_T_4; // @[ToAXI4.scala 200:45]
  assign queue_arw_deq_io_enq_bits_id = 7'h41 == auto_in_a_bits_source ? 7'h41 : _GEN_66; // @[ToAXI4.scala 169:{17,17}]
  assign queue_arw_deq_io_enq_bits_addr = auto_in_a_bits_address; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign queue_arw_deq_io_enq_bits_len = _out_arw_bits_len_T_3[13:6]; // @[ToAXI4.scala 171:84]
  assign queue_arw_deq_io_enq_bits_size = auto_in_a_bits_size >= 3'h6 ? 3'h6 : auto_in_a_bits_size; // @[ToAXI4.scala 172:23]
  assign queue_arw_deq_io_enq_bits_echo_tl_state_source = auto_in_a_bits_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign queue_arw_deq_io_enq_bits_wen = ~auto_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  assign queue_arw_deq_io_deq_ready = queue_arw_bits_wen ? auto_out_aw_ready : auto_out_ar_ready; // @[ToAXI4.scala 160:29]
  always @(posedge clock) begin
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_66 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_66 <= _count_T_262 - dec_65; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_65 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_65 <= _count_T_258 - dec_64; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_64 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_64 <= _count_T_254 - dec_63; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_63 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_63 <= _count_T_250 - dec_62; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_62 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_62 <= _count_T_246 - dec_61; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_61 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_61 <= _count_T_242 - dec_60; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_60 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_60 <= _count_T_238 - dec_59; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_59 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_59 <= _count_T_234 - dec_58; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_58 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_58 <= _count_T_230 - dec_57; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_57 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_57 <= _count_T_226 - dec_56; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_56 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_56 <= _count_T_222 - dec_55; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_55 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_55 <= _count_T_218 - dec_54; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_54 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_54 <= _count_T_214 - dec_53; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_53 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_53 <= _count_T_210 - dec_52; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_52 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_52 <= _count_T_206 - dec_51; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_51 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_51 <= _count_T_202 - dec_50; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_50 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_50 <= _count_T_198 - dec_49; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_49 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_49 <= _count_T_194 - dec_48; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_48 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_48 <= _count_T_190 - dec_47; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_47 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_47 <= _count_T_186 - dec_46; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_46 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_46 <= _count_T_182 - dec_45; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_45 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_45 <= _count_T_178 - dec_44; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_44 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_44 <= _count_T_174 - dec_43; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_43 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_43 <= _count_T_170 - dec_42; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_42 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_42 <= _count_T_166 - dec_41; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_41 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_41 <= _count_T_162 - dec_40; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_40 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_40 <= _count_T_158 - dec_39; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_39 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_39 <= _count_T_154 - dec_38; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_38 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_38 <= _count_T_150 - dec_37; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_37 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_37 <= _count_T_146 - dec_36; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_36 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_36 <= _count_T_142 - dec_35; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_35 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_35 <= _count_T_138 - dec_34; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_34 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_34 <= _count_T_134 - dec_33; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_33 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_33 <= _count_T_130 - dec_32; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_32 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_32 <= _count_T_126 - dec_31; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_31 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_31 <= _count_T_122 - dec_30; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_30 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_30 <= _count_T_118 - dec_29; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_29 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_29 <= _count_T_114 - dec_28; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_28 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_28 <= _count_T_110 - dec_27; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_27 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_27 <= _count_T_106 - dec_26; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_26 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_26 <= _count_T_102 - dec_25; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_25 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_25 <= _count_T_98 - dec_24; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_24 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_24 <= _count_T_94 - dec_23; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_23 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_23 <= _count_T_90 - dec_22; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_22 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_22 <= _count_T_86 - dec_21; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_21 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_21 <= _count_T_82 - dec_20; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_20 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_20 <= _count_T_78 - dec_19; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_19 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_19 <= _count_T_74 - dec_18; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_18 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_18 <= _count_T_70 - dec_17; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_17 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_17 <= _count_T_66 - dec_16; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_16 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_16 <= _count_T_62 - dec_15; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_15 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_15 <= _count_T_58 - dec_14; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_14 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_14 <= _count_T_54 - dec_13; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_13 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_13 <= _count_T_50 - dec_12; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_12 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_12 <= _count_T_46 - dec_11; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_11 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_11 <= _count_T_42 - dec_10; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_10 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_10 <= _count_T_38 - dec_9; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_9 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_9 <= _count_T_34 - dec_8; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_8 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_8 <= _count_T_30 - dec_7; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_7 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_7 <= _count_T_26 - dec_6; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_6 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_6 <= _count_T_22 - dec_5; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_5 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_5 <= _count_T_18 - dec_4; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_4 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_4 <= _count_T_14 - dec_3; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_3 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_3 <= _count_T_10 - dec_2; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_2 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_2 <= _count_T_6 - dec_1; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[ToAXI4.scala 257:28]
      count_1 <= 1'h0; // @[ToAXI4.scala 257:28]
    end else begin
      count_1 <= _count_T_2 - dec; // @[ToAXI4.scala 263:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      counter <= 1'h0; // @[Edges.scala 228:27]
    end else if (done) begin // @[Edges.scala 234:17]
      if (a_first) begin // @[Edges.scala 235:21]
        counter <= 1'h0;
      end else begin
        counter <= counter1;
      end
    end
    if (reset) begin // @[ToAXI4.scala 209:30]
      r_holds_d <= 1'h0; // @[ToAXI4.scala 209:30]
    end else if (_T_2) begin // @[ToAXI4.scala 210:27]
      r_holds_d <= ~auto_out_r_bits_last; // @[ToAXI4.scala 210:39]
    end
    if (auto_out_b_valid & ~x1_b_ready) begin // @[ToAXI4.scala 213:42]
      b_delay <= _b_delay_T_1; // @[ToAXI4.scala 214:17]
    end else begin
      b_delay <= 3'h0; // @[ToAXI4.scala 216:17]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec | count_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec | count_1) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc | idle)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc | idle) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_1 | count_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_1 | count_2) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_1 | idle_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_1 | idle_1) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_2 | count_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_2 | count_3) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_2 | idle_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_2 | idle_2) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_3 | count_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_3 | count_4) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_3 | idle_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_3 | idle_3) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_4 | count_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_4 | count_5) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_4 | idle_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_4 | idle_4) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_5 | count_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_5 | count_6) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_5 | idle_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_5 | idle_5) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_6 | count_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_6 | count_7) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_6 | idle_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_6 | idle_6) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_7 | count_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_7 | count_8) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_7 | idle_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_7 | idle_7) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_8 | count_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_8 | count_9) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_8 | idle_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_8 | idle_8) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_9 | count_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_9 | count_10) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_9 | idle_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_9 | idle_9) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_10 | count_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_10 | count_11) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_10 | idle_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_10 | idle_10) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_11 | count_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_11 | count_12) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_11 | idle_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_11 | idle_11) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_12 | count_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_12 | count_13) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_12 | idle_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_12 | idle_12) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_13 | count_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_13 | count_14) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_13 | idle_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_13 | idle_13) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_14 | count_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_14 | count_15) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_14 | idle_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_14 | idle_14) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_15 | count_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_15 | count_16) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_15 | idle_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_15 | idle_15) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_16 | count_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_16 | count_17) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_16 | idle_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_16 | idle_16) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_17 | count_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_17 | count_18) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_17 | idle_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_17 | idle_17) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_18 | count_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_18 | count_19) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_18 | idle_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_18 | idle_18) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_19 | count_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_19 | count_20) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_19 | idle_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_19 | idle_19) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_20 | count_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_20 | count_21) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_20 | idle_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_20 | idle_20) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_21 | count_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_21 | count_22) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_21 | idle_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_21 | idle_21) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_22 | count_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_22 | count_23) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_22 | idle_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_22 | idle_22) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_23 | count_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_23 | count_24) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_23 | idle_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_23 | idle_23) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_24 | count_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_24 | count_25) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_24 | idle_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_24 | idle_24) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_25 | count_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_25 | count_26) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_25 | idle_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_25 | idle_25) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_26 | count_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_26 | count_27) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_26 | idle_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_26 | idle_26) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_27 | count_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_27 | count_28) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_27 | idle_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_27 | idle_27) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_28 | count_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_28 | count_29) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_28 | idle_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_28 | idle_28) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_29 | count_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_29 | count_30) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_29 | idle_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_29 | idle_29) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_30 | count_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_30 | count_31) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_30 | idle_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_30 | idle_30) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_31 | count_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_31 | count_32) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_31 | idle_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_31 | idle_31) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_32 | count_33)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_32 | count_33) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_32 | idle_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_32 | idle_32) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_33 | count_34)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_33 | count_34) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_33 | idle_33)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_33 | idle_33) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_34 | count_35)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_34 | count_35) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_34 | idle_34)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_34 | idle_34) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_35 | count_36)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_35 | count_36) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_35 | idle_35)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_35 | idle_35) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_36 | count_37)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_36 | count_37) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_36 | idle_36)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_36 | idle_36) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_37 | count_38)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_37 | count_38) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_37 | idle_37)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_37 | idle_37) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_38 | count_39)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_38 | count_39) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_38 | idle_38)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_38 | idle_38) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_39 | count_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_39 | count_40) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_39 | idle_39)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_39 | idle_39) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_40 | count_41)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_40 | count_41) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_40 | idle_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_40 | idle_40) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_41 | count_42)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_41 | count_42) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_41 | idle_41)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_41 | idle_41) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_42 | count_43)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_42 | count_43) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_42 | idle_42)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_42 | idle_42) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_43 | count_44)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_43 | count_44) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_43 | idle_43)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_43 | idle_43) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_44 | count_45)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_44 | count_45) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_44 | idle_44)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_44 | idle_44) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_45 | count_46)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_45 | count_46) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_45 | idle_45)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_45 | idle_45) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_46 | count_47)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_46 | count_47) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_46 | idle_46)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_46 | idle_46) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_47 | count_48)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_47 | count_48) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_47 | idle_47)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_47 | idle_47) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_48 | count_49)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_48 | count_49) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_48 | idle_48)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_48 | idle_48) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_49 | count_50)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_49 | count_50) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_49 | idle_49)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_49 | idle_49) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_50 | count_51)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_50 | count_51) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_50 | idle_50)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_50 | idle_50) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_51 | count_52)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_51 | count_52) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_51 | idle_51)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_51 | idle_51) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_52 | count_53)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_52 | count_53) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_52 | idle_52)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_52 | idle_52) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_53 | count_54)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_53 | count_54) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_53 | idle_53)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_53 | idle_53) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_54 | count_55)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_54 | count_55) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_54 | idle_54)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_54 | idle_54) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_55 | count_56)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_55 | count_56) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_55 | idle_55)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_55 | idle_55) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_56 | count_57)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_56 | count_57) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_56 | idle_56)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_56 | idle_56) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_57 | count_58)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_57 | count_58) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_57 | idle_57)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_57 | idle_57) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_58 | count_59)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_58 | count_59) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_58 | idle_58)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_58 | idle_58) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_59 | count_60)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_59 | count_60) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_59 | idle_59)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_59 | idle_59) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_60 | count_61)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_60 | count_61) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_60 | idle_60)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_60 | idle_60) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_61 | count_62)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_61 | count_62) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_61 | idle_61)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_61 | idle_61) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_62 | count_63)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_62 | count_63) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_62 | idle_62)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_62 | idle_62) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_63 | count_64)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_63 | count_64) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_63 | idle_63)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_63 | idle_63) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_64 | count_65)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_64 | count_65) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_64 | idle_64)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_64 | idle_64) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_65 | count_66)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:265 assert (!dec || count =/= 0.U)        // underflow\n"); // @[ToAXI4.scala 265:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_65 | count_66) & ~reset) begin
          $fatal; // @[ToAXI4.scala 265:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_65 | idle_65)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:266 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[ToAXI4.scala 266:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_65 | idle_65) & _T_10) begin
          $fatal; // @[ToAXI4.scala 266:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_20(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [1:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [1:0] io_deq_bits
);
  reg [1:0] ram [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_12 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 318:26 280:27 318:35]
  wire  do_enq = empty ? _GEN_12 : _do_enq_T; // @[Decoupled.scala 315:17 280:27]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 315:17 317:14 281:27]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 302:16 314:{24,39}]
  assign io_deq_bits = empty ? io_enq_bits : ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      if (empty) begin // @[Decoupled.scala 315:17]
        if (io_deq_ready) begin // @[Decoupled.scala 318:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 318:35]
        end else begin
          maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
        end
      end else begin
        maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
      end
    end
  end
endmodule
module AXI4Xbar(
  input          clock,
  input          reset,
  output         auto_in_1_aw_ready,
  input          auto_in_1_aw_valid,
  input  [5:0]   auto_in_1_aw_bits_id,
  input  [33:0]  auto_in_1_aw_bits_addr,
  input  [7:0]   auto_in_1_aw_bits_len,
  input  [2:0]   auto_in_1_aw_bits_size,
  input  [1:0]   auto_in_1_aw_bits_burst,
  input          auto_in_1_aw_bits_lock,
  input  [3:0]   auto_in_1_aw_bits_cache,
  input  [2:0]   auto_in_1_aw_bits_prot,
  input  [3:0]   auto_in_1_aw_bits_qos,
  output         auto_in_1_w_ready,
  input          auto_in_1_w_valid,
  input  [511:0] auto_in_1_w_bits_data,
  input  [63:0]  auto_in_1_w_bits_strb,
  input          auto_in_1_w_bits_last,
  input          auto_in_1_b_ready,
  output         auto_in_1_b_valid,
  output [5:0]   auto_in_1_b_bits_id,
  output [1:0]   auto_in_1_b_bits_resp,
  output         auto_in_1_ar_ready,
  input          auto_in_1_ar_valid,
  input  [5:0]   auto_in_1_ar_bits_id,
  input  [33:0]  auto_in_1_ar_bits_addr,
  input  [7:0]   auto_in_1_ar_bits_len,
  input  [2:0]   auto_in_1_ar_bits_size,
  input  [1:0]   auto_in_1_ar_bits_burst,
  input          auto_in_1_ar_bits_lock,
  input  [3:0]   auto_in_1_ar_bits_cache,
  input  [2:0]   auto_in_1_ar_bits_prot,
  input  [3:0]   auto_in_1_ar_bits_qos,
  input          auto_in_1_r_ready,
  output         auto_in_1_r_valid,
  output [5:0]   auto_in_1_r_bits_id,
  output [511:0] auto_in_1_r_bits_data,
  output [1:0]   auto_in_1_r_bits_resp,
  output         auto_in_1_r_bits_last,
  output         auto_in_0_aw_ready,
  input          auto_in_0_aw_valid,
  input  [6:0]   auto_in_0_aw_bits_id,
  input  [33:0]  auto_in_0_aw_bits_addr,
  input  [7:0]   auto_in_0_aw_bits_len,
  input  [2:0]   auto_in_0_aw_bits_size,
  input  [1:0]   auto_in_0_aw_bits_burst,
  input          auto_in_0_aw_bits_lock,
  input  [3:0]   auto_in_0_aw_bits_cache,
  input  [2:0]   auto_in_0_aw_bits_prot,
  input  [3:0]   auto_in_0_aw_bits_qos,
  input  [6:0]   auto_in_0_aw_bits_echo_tl_state_source,
  output         auto_in_0_w_ready,
  input          auto_in_0_w_valid,
  input  [511:0] auto_in_0_w_bits_data,
  input  [63:0]  auto_in_0_w_bits_strb,
  input          auto_in_0_w_bits_last,
  input          auto_in_0_b_ready,
  output         auto_in_0_b_valid,
  output [6:0]   auto_in_0_b_bits_id,
  output [6:0]   auto_in_0_b_bits_echo_tl_state_source,
  output         auto_in_0_ar_ready,
  input          auto_in_0_ar_valid,
  input  [6:0]   auto_in_0_ar_bits_id,
  input  [33:0]  auto_in_0_ar_bits_addr,
  input  [7:0]   auto_in_0_ar_bits_len,
  input  [2:0]   auto_in_0_ar_bits_size,
  input  [1:0]   auto_in_0_ar_bits_burst,
  input          auto_in_0_ar_bits_lock,
  input  [3:0]   auto_in_0_ar_bits_cache,
  input  [2:0]   auto_in_0_ar_bits_prot,
  input  [3:0]   auto_in_0_ar_bits_qos,
  input  [6:0]   auto_in_0_ar_bits_echo_tl_state_source,
  input          auto_in_0_r_ready,
  output         auto_in_0_r_valid,
  output [6:0]   auto_in_0_r_bits_id,
  output [511:0] auto_in_0_r_bits_data,
  output [6:0]   auto_in_0_r_bits_echo_tl_state_source,
  output         auto_in_0_r_bits_last,
  input          auto_out_aw_ready,
  output         auto_out_aw_valid,
  output [7:0]   auto_out_aw_bits_id,
  output [33:0]  auto_out_aw_bits_addr,
  output [7:0]   auto_out_aw_bits_len,
  output [2:0]   auto_out_aw_bits_size,
  output [1:0]   auto_out_aw_bits_burst,
  output         auto_out_aw_bits_lock,
  output [3:0]   auto_out_aw_bits_cache,
  output [2:0]   auto_out_aw_bits_prot,
  output [3:0]   auto_out_aw_bits_qos,
  output [6:0]   auto_out_aw_bits_echo_tl_state_source,
  input          auto_out_w_ready,
  output         auto_out_w_valid,
  output [511:0] auto_out_w_bits_data,
  output [63:0]  auto_out_w_bits_strb,
  output         auto_out_w_bits_last,
  output         auto_out_b_ready,
  input          auto_out_b_valid,
  input  [7:0]   auto_out_b_bits_id,
  input  [1:0]   auto_out_b_bits_resp,
  input  [6:0]   auto_out_b_bits_echo_tl_state_source,
  input          auto_out_ar_ready,
  output         auto_out_ar_valid,
  output [7:0]   auto_out_ar_bits_id,
  output [33:0]  auto_out_ar_bits_addr,
  output [7:0]   auto_out_ar_bits_len,
  output [2:0]   auto_out_ar_bits_size,
  output [1:0]   auto_out_ar_bits_burst,
  output         auto_out_ar_bits_lock,
  output [3:0]   auto_out_ar_bits_cache,
  output [2:0]   auto_out_ar_bits_prot,
  output [3:0]   auto_out_ar_bits_qos,
  output [6:0]   auto_out_ar_bits_echo_tl_state_source,
  output         auto_out_r_ready,
  input          auto_out_r_valid,
  input  [7:0]   auto_out_r_bits_id,
  input  [511:0] auto_out_r_bits_data,
  input  [1:0]   auto_out_r_bits_resp,
  input  [6:0]   auto_out_r_bits_echo_tl_state_source,
  input          auto_out_r_bits_last
);
  wire  awOut_0_clock; // @[Xbar.scala 72:47]
  wire  awOut_0_reset; // @[Xbar.scala 72:47]
  wire  awOut_0_io_enq_ready; // @[Xbar.scala 72:47]
  wire  awOut_0_io_enq_valid; // @[Xbar.scala 72:47]
  wire [1:0] awOut_0_io_enq_bits; // @[Xbar.scala 72:47]
  wire  awOut_0_io_deq_ready; // @[Xbar.scala 72:47]
  wire  awOut_0_io_deq_valid; // @[Xbar.scala 72:47]
  wire [1:0] awOut_0_io_deq_bits; // @[Xbar.scala 72:47]
  wire  requestROI_0_0 = ~auto_out_r_bits_id[7]; // @[Parameters.scala 54:32]
  wire  requestROI_0_1 = auto_out_r_bits_id[7:6] == 2'h2; // @[Parameters.scala 54:32]
  wire  requestBOI_0_0 = ~auto_out_b_bits_id[7]; // @[Parameters.scala 54:32]
  wire  requestBOI_0_1 = auto_out_b_bits_id[7:6] == 2'h2; // @[Parameters.scala 54:32]
  wire [7:0] _GEN_16 = {{2'd0}, auto_in_1_aw_bits_id}; // @[Xbar.scala 95:47]
  wire [7:0] in_1_aw_bits_id = _GEN_16 | 8'h80; // @[Xbar.scala 95:47]
  wire [7:0] _GEN_17 = {{2'd0}, auto_in_1_ar_bits_id}; // @[Xbar.scala 96:47]
  wire [7:0] in_1_ar_bits_id = _GEN_17 | 8'h80; // @[Xbar.scala 96:47]
  reg  latched; // @[Xbar.scala 176:30]
  wire  _x1_aw_valid_T = latched | awOut_0_io_enq_ready; // @[Xbar.scala 177:59]
  reg  awOut_0_io_enq_bits_idle; // @[Xbar.scala 262:23]
  wire  awOut_0_io_enq_bits_anyValid = auto_in_0_aw_valid | auto_in_1_aw_valid; // @[Xbar.scala 266:36]
  reg  awOut_0_io_enq_bits_state_0; // @[Xbar.scala 281:24]
  reg  awOut_0_io_enq_bits_state_1; // @[Xbar.scala 281:24]
  wire  _awOut_0_io_enq_bits_out_0_aw_valid_T_2 = awOut_0_io_enq_bits_state_0 & auto_in_0_aw_valid |
    awOut_0_io_enq_bits_state_1 & auto_in_1_aw_valid; // @[Mux.scala 27:73]
  wire  out_0_aw_valid = awOut_0_io_enq_bits_idle ? awOut_0_io_enq_bits_anyValid :
    _awOut_0_io_enq_bits_out_0_aw_valid_T_2; // @[Xbar.scala 298:22]
  wire  out_0_aw_ready = auto_out_aw_ready & _x1_aw_valid_T; // @[Xbar.scala 178:47]
  wire  _T = awOut_0_io_enq_ready & awOut_0_io_enq_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_0 = _T | latched; // @[Xbar.scala 176:30 180:{37,47}]
  wire  _T_1 = out_0_aw_ready & out_0_aw_valid; // @[Decoupled.scala 51:35]
  wire  out_0_w_valid = awOut_0_io_deq_bits[0] & auto_in_0_w_valid | awOut_0_io_deq_bits[1] & auto_in_1_w_valid; // @[Mux.scala 27:73]
  wire  out_0_w_ready = auto_out_w_ready & awOut_0_io_deq_valid; // @[Xbar.scala 185:45]
  wire  out_0_w_bits_last = awOut_0_io_deq_bits[0] & auto_in_0_w_bits_last | awOut_0_io_deq_bits[1] &
    auto_in_1_w_bits_last; // @[Mux.scala 27:73]
  wire  portsRIO_filtered_0_valid = auto_out_r_valid & requestROI_0_0; // @[Xbar.scala 242:40]
  wire  portsRIO_filtered_1_valid = auto_out_r_valid & requestROI_0_1; // @[Xbar.scala 242:40]
  wire  portsBIO_filtered_0_valid = auto_out_b_valid & requestBOI_0_0; // @[Xbar.scala 242:40]
  wire  portsBIO_filtered_1_valid = auto_out_b_valid & requestBOI_0_1; // @[Xbar.scala 242:40]
  wire [1:0] awOut_0_io_enq_bits_readys_valid = {auto_in_1_aw_valid,auto_in_0_aw_valid}; // @[Cat.scala 33:92]
  wire  _awOut_0_io_enq_bits_readys_T_3 = ~reset; // @[Arbiter.scala 23:12]
  reg [1:0] awOut_0_io_enq_bits_readys_mask; // @[Arbiter.scala 24:23]
  wire [1:0] _awOut_0_io_enq_bits_readys_filter_T = ~awOut_0_io_enq_bits_readys_mask; // @[Arbiter.scala 25:30]
  wire [1:0] _awOut_0_io_enq_bits_readys_filter_T_1 = awOut_0_io_enq_bits_readys_valid &
    _awOut_0_io_enq_bits_readys_filter_T; // @[Arbiter.scala 25:28]
  wire [3:0] awOut_0_io_enq_bits_readys_filter = {_awOut_0_io_enq_bits_readys_filter_T_1,auto_in_1_aw_valid,
    auto_in_0_aw_valid}; // @[Cat.scala 33:92]
  wire [3:0] _GEN_18 = {{1'd0}, awOut_0_io_enq_bits_readys_filter[3:1]}; // @[package.scala 254:43]
  wire [3:0] _awOut_0_io_enq_bits_readys_unready_T_1 = awOut_0_io_enq_bits_readys_filter | _GEN_18; // @[package.scala 254:43]
  wire [3:0] _awOut_0_io_enq_bits_readys_unready_T_4 = {awOut_0_io_enq_bits_readys_mask, 2'h0}; // @[Arbiter.scala 26:66]
  wire [3:0] _GEN_19 = {{1'd0}, _awOut_0_io_enq_bits_readys_unready_T_1[3:1]}; // @[Arbiter.scala 26:58]
  wire [3:0] awOut_0_io_enq_bits_readys_unready = _GEN_19 | _awOut_0_io_enq_bits_readys_unready_T_4; // @[Arbiter.scala 26:58]
  wire [1:0] _awOut_0_io_enq_bits_readys_readys_T_2 = awOut_0_io_enq_bits_readys_unready[3:2] &
    awOut_0_io_enq_bits_readys_unready[1:0]; // @[Arbiter.scala 27:39]
  wire [1:0] awOut_0_io_enq_bits_readys_readys = ~_awOut_0_io_enq_bits_readys_readys_T_2; // @[Arbiter.scala 27:18]
  wire [1:0] _awOut_0_io_enq_bits_readys_mask_T = awOut_0_io_enq_bits_readys_readys & awOut_0_io_enq_bits_readys_valid; // @[Arbiter.scala 29:29]
  wire [2:0] _awOut_0_io_enq_bits_readys_mask_T_1 = {_awOut_0_io_enq_bits_readys_mask_T, 1'h0}; // @[package.scala 245:48]
  wire [1:0] _awOut_0_io_enq_bits_readys_mask_T_3 = _awOut_0_io_enq_bits_readys_mask_T |
    _awOut_0_io_enq_bits_readys_mask_T_1[1:0]; // @[package.scala 245:43]
  wire  awOut_0_io_enq_bits_readys_0 = awOut_0_io_enq_bits_readys_readys[0]; // @[Xbar.scala 268:73]
  wire  awOut_0_io_enq_bits_readys_1 = awOut_0_io_enq_bits_readys_readys[1]; // @[Xbar.scala 268:73]
  wire  awOut_0_io_enq_bits_winner_0 = awOut_0_io_enq_bits_readys_0 & auto_in_0_aw_valid; // @[Xbar.scala 270:67]
  wire  awOut_0_io_enq_bits_winner_1 = awOut_0_io_enq_bits_readys_1 & auto_in_1_aw_valid; // @[Xbar.scala 270:67]
  wire  _awOut_0_io_enq_bits_prefixOR_T = awOut_0_io_enq_bits_winner_0 | awOut_0_io_enq_bits_winner_1; // @[Xbar.scala 275:46]
  wire  awOut_0_io_enq_bits_muxState_0 = awOut_0_io_enq_bits_idle ? awOut_0_io_enq_bits_winner_0 :
    awOut_0_io_enq_bits_state_0; // @[Xbar.scala 282:23]
  wire  awOut_0_io_enq_bits_muxState_1 = awOut_0_io_enq_bits_idle ? awOut_0_io_enq_bits_winner_1 :
    awOut_0_io_enq_bits_state_1; // @[Xbar.scala 282:23]
  wire  _GEN_3 = awOut_0_io_enq_bits_anyValid ? 1'h0 : awOut_0_io_enq_bits_idle; // @[Xbar.scala 286:21 262:23 286:28]
  wire  _GEN_4 = _T_1 | _GEN_3; // @[Xbar.scala 287:{22,29}]
  wire  awOut_0_io_enq_bits_allowed_0 = awOut_0_io_enq_bits_idle ? awOut_0_io_enq_bits_readys_0 :
    awOut_0_io_enq_bits_state_0; // @[Xbar.scala 290:24]
  wire  awOut_0_io_enq_bits_allowed_1 = awOut_0_io_enq_bits_idle ? awOut_0_io_enq_bits_readys_1 :
    awOut_0_io_enq_bits_state_1; // @[Xbar.scala 290:24]
  wire [3:0] _awOut_0_io_enq_bits_T_23 = awOut_0_io_enq_bits_muxState_0 ? auto_in_0_aw_bits_qos : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _awOut_0_io_enq_bits_T_24 = awOut_0_io_enq_bits_muxState_1 ? auto_in_1_aw_bits_qos : 4'h0; // @[Mux.scala 27:73]
  wire [2:0] _awOut_0_io_enq_bits_T_26 = awOut_0_io_enq_bits_muxState_0 ? auto_in_0_aw_bits_prot : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _awOut_0_io_enq_bits_T_27 = awOut_0_io_enq_bits_muxState_1 ? auto_in_1_aw_bits_prot : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _awOut_0_io_enq_bits_T_29 = awOut_0_io_enq_bits_muxState_0 ? auto_in_0_aw_bits_cache : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _awOut_0_io_enq_bits_T_30 = awOut_0_io_enq_bits_muxState_1 ? auto_in_1_aw_bits_cache : 4'h0; // @[Mux.scala 27:73]
  wire [1:0] _awOut_0_io_enq_bits_T_35 = awOut_0_io_enq_bits_muxState_0 ? auto_in_0_aw_bits_burst : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _awOut_0_io_enq_bits_T_36 = awOut_0_io_enq_bits_muxState_1 ? auto_in_1_aw_bits_burst : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _awOut_0_io_enq_bits_T_38 = awOut_0_io_enq_bits_muxState_0 ? auto_in_0_aw_bits_size : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _awOut_0_io_enq_bits_T_39 = awOut_0_io_enq_bits_muxState_1 ? auto_in_1_aw_bits_size : 3'h0; // @[Mux.scala 27:73]
  wire [7:0] _awOut_0_io_enq_bits_T_41 = awOut_0_io_enq_bits_muxState_0 ? auto_in_0_aw_bits_len : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _awOut_0_io_enq_bits_T_42 = awOut_0_io_enq_bits_muxState_1 ? auto_in_1_aw_bits_len : 8'h0; // @[Mux.scala 27:73]
  wire [33:0] _awOut_0_io_enq_bits_T_44 = awOut_0_io_enq_bits_muxState_0 ? auto_in_0_aw_bits_addr : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _awOut_0_io_enq_bits_T_45 = awOut_0_io_enq_bits_muxState_1 ? auto_in_1_aw_bits_addr : 34'h0; // @[Mux.scala 27:73]
  wire [7:0] in_0_aw_bits_id = {{1'd0}, auto_in_0_aw_bits_id}; // @[Xbar.scala 87:18 95:24]
  wire [7:0] _awOut_0_io_enq_bits_T_47 = awOut_0_io_enq_bits_muxState_0 ? in_0_aw_bits_id : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _awOut_0_io_enq_bits_T_48 = awOut_0_io_enq_bits_muxState_1 ? in_1_aw_bits_id : 8'h0; // @[Mux.scala 27:73]
  reg  idle; // @[Xbar.scala 262:23]
  wire  anyValid = auto_in_0_ar_valid | auto_in_1_ar_valid; // @[Xbar.scala 266:36]
  wire [1:0] readys_valid = {auto_in_1_ar_valid,auto_in_0_ar_valid}; // @[Cat.scala 33:92]
  reg [1:0] readys_mask; // @[Arbiter.scala 24:23]
  wire [1:0] _readys_filter_T = ~readys_mask; // @[Arbiter.scala 25:30]
  wire [1:0] _readys_filter_T_1 = readys_valid & _readys_filter_T; // @[Arbiter.scala 25:28]
  wire [3:0] readys_filter = {_readys_filter_T_1,auto_in_1_ar_valid,auto_in_0_ar_valid}; // @[Cat.scala 33:92]
  wire [3:0] _GEN_20 = {{1'd0}, readys_filter[3:1]}; // @[package.scala 254:43]
  wire [3:0] _readys_unready_T_1 = readys_filter | _GEN_20; // @[package.scala 254:43]
  wire [3:0] _readys_unready_T_4 = {readys_mask, 2'h0}; // @[Arbiter.scala 26:66]
  wire [3:0] _GEN_21 = {{1'd0}, _readys_unready_T_1[3:1]}; // @[Arbiter.scala 26:58]
  wire [3:0] readys_unready = _GEN_21 | _readys_unready_T_4; // @[Arbiter.scala 26:58]
  wire [1:0] _readys_readys_T_2 = readys_unready[3:2] & readys_unready[1:0]; // @[Arbiter.scala 27:39]
  wire [1:0] readys_readys = ~_readys_readys_T_2; // @[Arbiter.scala 27:18]
  wire [1:0] _readys_mask_T = readys_readys & readys_valid; // @[Arbiter.scala 29:29]
  wire [2:0] _readys_mask_T_1 = {_readys_mask_T, 1'h0}; // @[package.scala 245:48]
  wire [1:0] _readys_mask_T_3 = _readys_mask_T | _readys_mask_T_1[1:0]; // @[package.scala 245:43]
  wire  readys__0 = readys_readys[0]; // @[Xbar.scala 268:73]
  wire  readys__1 = readys_readys[1]; // @[Xbar.scala 268:73]
  wire  winner__0 = readys__0 & auto_in_0_ar_valid; // @[Xbar.scala 270:67]
  wire  winner__1 = readys__1 & auto_in_1_ar_valid; // @[Xbar.scala 270:67]
  wire  _prefixOR_T = winner__0 | winner__1; // @[Xbar.scala 275:46]
  reg  state__0; // @[Xbar.scala 281:24]
  reg  state__1; // @[Xbar.scala 281:24]
  wire  muxState__0 = idle ? winner__0 : state__0; // @[Xbar.scala 282:23]
  wire  muxState__1 = idle ? winner__1 : state__1; // @[Xbar.scala 282:23]
  wire  _GEN_6 = anyValid ? 1'h0 : idle; // @[Xbar.scala 286:21 262:23 286:28]
  wire  _out_0_ar_valid_T_2 = state__0 & auto_in_0_ar_valid | state__1 & auto_in_1_ar_valid; // @[Mux.scala 27:73]
  wire  out_0_ar_valid = idle ? anyValid : _out_0_ar_valid_T_2; // @[Xbar.scala 298:22]
  wire  _T_18 = auto_out_ar_ready & out_0_ar_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_7 = _T_18 | _GEN_6; // @[Xbar.scala 287:{22,29}]
  wire  allowed_0 = idle ? readys__0 : state__0; // @[Xbar.scala 290:24]
  wire  allowed_1 = idle ? readys__1 : state__1; // @[Xbar.scala 290:24]
  wire [3:0] _T_25 = muxState__0 ? auto_in_0_ar_bits_qos : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_26 = muxState__1 ? auto_in_1_ar_bits_qos : 4'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_28 = muxState__0 ? auto_in_0_ar_bits_prot : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_29 = muxState__1 ? auto_in_1_ar_bits_prot : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_31 = muxState__0 ? auto_in_0_ar_bits_cache : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_32 = muxState__1 ? auto_in_1_ar_bits_cache : 4'h0; // @[Mux.scala 27:73]
  wire [1:0] _T_37 = muxState__0 ? auto_in_0_ar_bits_burst : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _T_38 = muxState__1 ? auto_in_1_ar_bits_burst : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_40 = muxState__0 ? auto_in_0_ar_bits_size : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_41 = muxState__1 ? auto_in_1_ar_bits_size : 3'h0; // @[Mux.scala 27:73]
  wire [7:0] _T_43 = muxState__0 ? auto_in_0_ar_bits_len : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _T_44 = muxState__1 ? auto_in_1_ar_bits_len : 8'h0; // @[Mux.scala 27:73]
  wire [33:0] _T_46 = muxState__0 ? auto_in_0_ar_bits_addr : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _T_47 = muxState__1 ? auto_in_1_ar_bits_addr : 34'h0; // @[Mux.scala 27:73]
  wire [7:0] in_0_ar_bits_id = {{1'd0}, auto_in_0_ar_bits_id}; // @[Xbar.scala 87:18 96:24]
  wire [7:0] _T_49 = muxState__0 ? in_0_ar_bits_id : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _T_50 = muxState__1 ? in_1_ar_bits_id : 8'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_57 = awOut_0_io_deq_bits[0] ? auto_in_0_w_bits_strb : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_58 = awOut_0_io_deq_bits[1] ? auto_in_1_w_bits_strb : 64'h0; // @[Mux.scala 27:73]
  wire [511:0] _T_60 = awOut_0_io_deq_bits[0] ? auto_in_0_w_bits_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _T_61 = awOut_0_io_deq_bits[1] ? auto_in_1_w_bits_data : 512'h0; // @[Mux.scala 27:73]
  wire  _T_64 = ~portsRIO_filtered_0_valid; // @[Xbar.scala 276:60]
  wire  _T_76 = ~portsBIO_filtered_0_valid; // @[Xbar.scala 276:60]
  wire  _T_88 = ~portsRIO_filtered_1_valid; // @[Xbar.scala 276:60]
  wire  _T_100 = ~portsBIO_filtered_1_valid; // @[Xbar.scala 276:60]
  Queue_20 awOut_0 ( // @[Xbar.scala 72:47]
    .clock(awOut_0_clock),
    .reset(awOut_0_reset),
    .io_enq_ready(awOut_0_io_enq_ready),
    .io_enq_valid(awOut_0_io_enq_valid),
    .io_enq_bits(awOut_0_io_enq_bits),
    .io_deq_ready(awOut_0_io_deq_ready),
    .io_deq_valid(awOut_0_io_deq_valid),
    .io_deq_bits(awOut_0_io_deq_bits)
  );
  assign auto_in_1_aw_ready = out_0_aw_ready & awOut_0_io_enq_bits_allowed_1; // @[Xbar.scala 292:31]
  assign auto_in_1_w_ready = out_0_w_ready & awOut_0_io_deq_bits[1]; // @[Xbar.scala 210:37]
  assign auto_in_1_b_valid = auto_out_b_valid & requestBOI_0_1; // @[Xbar.scala 242:40]
  assign auto_in_1_b_bits_id = auto_out_b_bits_id[5:0]; // @[Xbar.scala 92:65]
  assign auto_in_1_b_bits_resp = auto_out_b_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_1_ar_ready = auto_out_ar_ready & allowed_1; // @[Xbar.scala 292:31]
  assign auto_in_1_r_valid = auto_out_r_valid & requestROI_0_1; // @[Xbar.scala 242:40]
  assign auto_in_1_r_bits_id = auto_out_r_bits_id[5:0]; // @[Xbar.scala 92:65]
  assign auto_in_1_r_bits_data = auto_out_r_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_1_r_bits_resp = auto_out_r_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_1_r_bits_last = auto_out_r_bits_last; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_0_aw_ready = out_0_aw_ready & awOut_0_io_enq_bits_allowed_0; // @[Xbar.scala 292:31]
  assign auto_in_0_w_ready = out_0_w_ready & awOut_0_io_deq_bits[0]; // @[Xbar.scala 210:37]
  assign auto_in_0_b_valid = auto_out_b_valid & requestBOI_0_0; // @[Xbar.scala 242:40]
  assign auto_in_0_b_bits_id = auto_out_b_bits_id[6:0]; // @[Xbar.scala 92:65]
  assign auto_in_0_b_bits_echo_tl_state_source = auto_out_b_bits_echo_tl_state_source; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_0_ar_ready = auto_out_ar_ready & allowed_0; // @[Xbar.scala 292:31]
  assign auto_in_0_r_valid = auto_out_r_valid & requestROI_0_0; // @[Xbar.scala 242:40]
  assign auto_in_0_r_bits_id = auto_out_r_bits_id[6:0]; // @[Xbar.scala 92:65]
  assign auto_in_0_r_bits_data = auto_out_r_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_0_r_bits_echo_tl_state_source = auto_out_r_bits_echo_tl_state_source; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_0_r_bits_last = auto_out_r_bits_last; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_out_aw_valid = out_0_aw_valid & (latched | awOut_0_io_enq_ready); // @[Xbar.scala 177:47]
  assign auto_out_aw_bits_id = _awOut_0_io_enq_bits_T_47 | _awOut_0_io_enq_bits_T_48; // @[Mux.scala 27:73]
  assign auto_out_aw_bits_addr = _awOut_0_io_enq_bits_T_44 | _awOut_0_io_enq_bits_T_45; // @[Mux.scala 27:73]
  assign auto_out_aw_bits_len = _awOut_0_io_enq_bits_T_41 | _awOut_0_io_enq_bits_T_42; // @[Mux.scala 27:73]
  assign auto_out_aw_bits_size = _awOut_0_io_enq_bits_T_38 | _awOut_0_io_enq_bits_T_39; // @[Mux.scala 27:73]
  assign auto_out_aw_bits_burst = _awOut_0_io_enq_bits_T_35 | _awOut_0_io_enq_bits_T_36; // @[Mux.scala 27:73]
  assign auto_out_aw_bits_lock = awOut_0_io_enq_bits_muxState_0 & auto_in_0_aw_bits_lock |
    awOut_0_io_enq_bits_muxState_1 & auto_in_1_aw_bits_lock; // @[Mux.scala 27:73]
  assign auto_out_aw_bits_cache = _awOut_0_io_enq_bits_T_29 | _awOut_0_io_enq_bits_T_30; // @[Mux.scala 27:73]
  assign auto_out_aw_bits_prot = _awOut_0_io_enq_bits_T_26 | _awOut_0_io_enq_bits_T_27; // @[Mux.scala 27:73]
  assign auto_out_aw_bits_qos = _awOut_0_io_enq_bits_T_23 | _awOut_0_io_enq_bits_T_24; // @[Mux.scala 27:73]
  assign auto_out_aw_bits_echo_tl_state_source = awOut_0_io_enq_bits_muxState_0 ? auto_in_0_aw_bits_echo_tl_state_source
     : 7'h0; // @[Mux.scala 27:73]
  assign auto_out_w_valid = out_0_w_valid & awOut_0_io_deq_valid; // @[Xbar.scala 184:45]
  assign auto_out_w_bits_data = _T_60 | _T_61; // @[Mux.scala 27:73]
  assign auto_out_w_bits_strb = _T_57 | _T_58; // @[Mux.scala 27:73]
  assign auto_out_w_bits_last = awOut_0_io_deq_bits[0] & auto_in_0_w_bits_last | awOut_0_io_deq_bits[1] &
    auto_in_1_w_bits_last; // @[Mux.scala 27:73]
  assign auto_out_b_ready = requestBOI_0_0 & auto_in_0_b_ready | requestBOI_0_1 & auto_in_1_b_ready; // @[Mux.scala 27:73]
  assign auto_out_ar_valid = idle ? anyValid : _out_0_ar_valid_T_2; // @[Xbar.scala 298:22]
  assign auto_out_ar_bits_id = _T_49 | _T_50; // @[Mux.scala 27:73]
  assign auto_out_ar_bits_addr = _T_46 | _T_47; // @[Mux.scala 27:73]
  assign auto_out_ar_bits_len = _T_43 | _T_44; // @[Mux.scala 27:73]
  assign auto_out_ar_bits_size = _T_40 | _T_41; // @[Mux.scala 27:73]
  assign auto_out_ar_bits_burst = _T_37 | _T_38; // @[Mux.scala 27:73]
  assign auto_out_ar_bits_lock = muxState__0 & auto_in_0_ar_bits_lock | muxState__1 & auto_in_1_ar_bits_lock; // @[Mux.scala 27:73]
  assign auto_out_ar_bits_cache = _T_31 | _T_32; // @[Mux.scala 27:73]
  assign auto_out_ar_bits_prot = _T_28 | _T_29; // @[Mux.scala 27:73]
  assign auto_out_ar_bits_qos = _T_25 | _T_26; // @[Mux.scala 27:73]
  assign auto_out_ar_bits_echo_tl_state_source = muxState__0 ? auto_in_0_ar_bits_echo_tl_state_source : 7'h0; // @[Mux.scala 27:73]
  assign auto_out_r_ready = requestROI_0_0 & auto_in_0_r_ready | requestROI_0_1 & auto_in_1_r_ready; // @[Mux.scala 27:73]
  assign awOut_0_clock = clock;
  assign awOut_0_reset = reset;
  assign awOut_0_io_enq_valid = out_0_aw_valid & ~latched; // @[Xbar.scala 179:50]
  assign awOut_0_io_enq_bits = {awOut_0_io_enq_bits_muxState_1,awOut_0_io_enq_bits_muxState_0}; // @[Xbar.scala 203:81]
  assign awOut_0_io_deq_ready = out_0_w_valid & out_0_w_bits_last & auto_out_w_ready; // @[Xbar.scala 186:71]
  always @(posedge clock) begin
    if (reset) begin // @[Xbar.scala 176:30]
      latched <= 1'h0; // @[Xbar.scala 176:30]
    end else if (_T_1) begin // @[Xbar.scala 181:31]
      latched <= 1'h0; // @[Xbar.scala 181:41]
    end else begin
      latched <= _GEN_0;
    end
    awOut_0_io_enq_bits_idle <= reset | _GEN_4; // @[Xbar.scala 262:{23,23}]
    if (reset) begin // @[Xbar.scala 281:24]
      awOut_0_io_enq_bits_state_0 <= 1'h0; // @[Xbar.scala 281:24]
    end else if (awOut_0_io_enq_bits_idle) begin // @[Xbar.scala 282:23]
      awOut_0_io_enq_bits_state_0 <= awOut_0_io_enq_bits_winner_0;
    end
    if (reset) begin // @[Xbar.scala 281:24]
      awOut_0_io_enq_bits_state_1 <= 1'h0; // @[Xbar.scala 281:24]
    end else if (awOut_0_io_enq_bits_idle) begin // @[Xbar.scala 282:23]
      awOut_0_io_enq_bits_state_1 <= awOut_0_io_enq_bits_winner_1;
    end
    if (reset) begin // @[Arbiter.scala 24:23]
      awOut_0_io_enq_bits_readys_mask <= 2'h3; // @[Arbiter.scala 24:23]
    end else if (awOut_0_io_enq_bits_idle & |awOut_0_io_enq_bits_readys_valid) begin // @[Arbiter.scala 28:32]
      awOut_0_io_enq_bits_readys_mask <= _awOut_0_io_enq_bits_readys_mask_T_3; // @[Arbiter.scala 29:12]
    end
    idle <= reset | _GEN_7; // @[Xbar.scala 262:{23,23}]
    if (reset) begin // @[Arbiter.scala 24:23]
      readys_mask <= 2'h3; // @[Arbiter.scala 24:23]
    end else if (idle & |readys_valid) begin // @[Arbiter.scala 28:32]
      readys_mask <= _readys_mask_T_3; // @[Arbiter.scala 29:12]
    end
    if (reset) begin // @[Xbar.scala 281:24]
      state__0 <= 1'h0; // @[Xbar.scala 281:24]
    end else if (idle) begin // @[Xbar.scala 282:23]
      state__0 <= winner__0;
    end
    if (reset) begin // @[Xbar.scala 281:24]
      state__1 <= 1'h0; // @[Xbar.scala 281:24]
    end else if (idle) begin // @[Xbar.scala 282:23]
      state__1 <= winner__1;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_awOut_0_io_enq_bits_readys_T_3 & ~(~awOut_0_io_enq_bits_winner_0 | ~awOut_0_io_enq_bits_winner_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Xbar.scala:276 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[Xbar.scala 276:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~awOut_0_io_enq_bits_winner_0 | ~awOut_0_io_enq_bits_winner_1) & _awOut_0_io_enq_bits_readys_T_3) begin
          $fatal; // @[Xbar.scala 276:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_awOut_0_io_enq_bits_readys_T_3 & ~(~awOut_0_io_enq_bits_anyValid | _awOut_0_io_enq_bits_prefixOR_T)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:278 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 278:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~awOut_0_io_enq_bits_anyValid | _awOut_0_io_enq_bits_prefixOR_T) & _awOut_0_io_enq_bits_readys_T_3) begin
          $fatal; // @[Xbar.scala 278:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_awOut_0_io_enq_bits_readys_T_3 & ~(~winner__0 | ~winner__1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Xbar.scala:276 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[Xbar.scala 276:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~winner__0 | ~winner__1) & _awOut_0_io_enq_bits_readys_T_3) begin
          $fatal; // @[Xbar.scala 276:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_awOut_0_io_enq_bits_readys_T_3 & ~(~anyValid | _prefixOR_T)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:278 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 278:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~anyValid | _prefixOR_T) & _awOut_0_io_enq_bits_readys_T_3) begin
          $fatal; // @[Xbar.scala 278:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_awOut_0_io_enq_bits_readys_T_3 & ~(_T_64 | portsRIO_filtered_0_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:278 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 278:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_64 | portsRIO_filtered_0_valid) & _awOut_0_io_enq_bits_readys_T_3) begin
          $fatal; // @[Xbar.scala 278:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_awOut_0_io_enq_bits_readys_T_3 & ~(_T_76 | portsBIO_filtered_0_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:278 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 278:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_76 | portsBIO_filtered_0_valid) & _awOut_0_io_enq_bits_readys_T_3) begin
          $fatal; // @[Xbar.scala 278:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_awOut_0_io_enq_bits_readys_T_3 & ~(_T_88 | portsRIO_filtered_1_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:278 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 278:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_88 | portsRIO_filtered_1_valid) & _awOut_0_io_enq_bits_readys_T_3) begin
          $fatal; // @[Xbar.scala 278:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_awOut_0_io_enq_bits_readys_T_3 & ~(_T_100 | portsBIO_filtered_1_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:278 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 278:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_100 | portsBIO_filtered_1_valid) & _awOut_0_io_enq_bits_readys_T_3) begin
          $fatal; // @[Xbar.scala 278:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module AXI4Xbar_1(
  input          clock,
  input          reset,
  output         auto_in_aw_ready,
  input          auto_in_aw_valid,
  input  [5:0]   auto_in_aw_bits_id,
  input  [33:0]  auto_in_aw_bits_addr,
  input  [7:0]   auto_in_aw_bits_len,
  input  [2:0]   auto_in_aw_bits_size,
  input  [1:0]   auto_in_aw_bits_burst,
  input          auto_in_aw_bits_lock,
  input  [3:0]   auto_in_aw_bits_cache,
  input  [2:0]   auto_in_aw_bits_prot,
  input  [3:0]   auto_in_aw_bits_qos,
  output         auto_in_w_ready,
  input          auto_in_w_valid,
  input  [511:0] auto_in_w_bits_data,
  input  [63:0]  auto_in_w_bits_strb,
  input          auto_in_w_bits_last,
  input          auto_in_b_ready,
  output         auto_in_b_valid,
  output [5:0]   auto_in_b_bits_id,
  output [1:0]   auto_in_b_bits_resp,
  output         auto_in_ar_ready,
  input          auto_in_ar_valid,
  input  [5:0]   auto_in_ar_bits_id,
  input  [33:0]  auto_in_ar_bits_addr,
  input  [7:0]   auto_in_ar_bits_len,
  input  [2:0]   auto_in_ar_bits_size,
  input  [1:0]   auto_in_ar_bits_burst,
  input          auto_in_ar_bits_lock,
  input  [3:0]   auto_in_ar_bits_cache,
  input  [2:0]   auto_in_ar_bits_prot,
  input  [3:0]   auto_in_ar_bits_qos,
  input          auto_in_r_ready,
  output         auto_in_r_valid,
  output [5:0]   auto_in_r_bits_id,
  output [511:0] auto_in_r_bits_data,
  output [1:0]   auto_in_r_bits_resp,
  output         auto_in_r_bits_last,
  input          auto_out_aw_ready,
  output         auto_out_aw_valid,
  output [5:0]   auto_out_aw_bits_id,
  output [33:0]  auto_out_aw_bits_addr,
  output [7:0]   auto_out_aw_bits_len,
  output [2:0]   auto_out_aw_bits_size,
  output [1:0]   auto_out_aw_bits_burst,
  output         auto_out_aw_bits_lock,
  output [3:0]   auto_out_aw_bits_cache,
  output [2:0]   auto_out_aw_bits_prot,
  output [3:0]   auto_out_aw_bits_qos,
  input          auto_out_w_ready,
  output         auto_out_w_valid,
  output [511:0] auto_out_w_bits_data,
  output [63:0]  auto_out_w_bits_strb,
  output         auto_out_w_bits_last,
  output         auto_out_b_ready,
  input          auto_out_b_valid,
  input  [5:0]   auto_out_b_bits_id,
  input  [1:0]   auto_out_b_bits_resp,
  input          auto_out_ar_ready,
  output         auto_out_ar_valid,
  output [5:0]   auto_out_ar_bits_id,
  output [33:0]  auto_out_ar_bits_addr,
  output [7:0]   auto_out_ar_bits_len,
  output [2:0]   auto_out_ar_bits_size,
  output [1:0]   auto_out_ar_bits_burst,
  output         auto_out_ar_bits_lock,
  output [3:0]   auto_out_ar_bits_cache,
  output [2:0]   auto_out_ar_bits_prot,
  output [3:0]   auto_out_ar_bits_qos,
  output         auto_out_r_ready,
  input          auto_out_r_valid,
  input  [5:0]   auto_out_r_bits_id,
  input  [511:0] auto_out_r_bits_data,
  input  [1:0]   auto_out_r_bits_resp,
  input          auto_out_r_bits_last
);
  wire  _awOut_0_io_enq_bits_T_1 = ~auto_in_aw_valid; // @[Xbar.scala 276:60]
  wire  _awOut_0_io_enq_bits_T_4 = ~reset; // @[Xbar.scala 276:11]
  wire  _T_1 = ~auto_in_ar_valid; // @[Xbar.scala 276:60]
  wire  _T_14 = ~auto_out_r_valid; // @[Xbar.scala 276:60]
  wire  _T_26 = ~auto_out_b_valid; // @[Xbar.scala 276:60]
  assign auto_in_aw_ready = auto_out_aw_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_w_ready = auto_out_w_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_b_valid = auto_out_b_valid; // @[Xbar.scala 298:22]
  assign auto_in_b_bits_id = auto_out_b_bits_id; // @[Xbar.scala 92:65]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_ar_ready = auto_out_ar_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_valid = auto_out_r_valid; // @[Xbar.scala 298:22]
  assign auto_in_r_bits_id = auto_out_r_bits_id; // @[Xbar.scala 92:65]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_bits_last = auto_out_r_bits_last; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_out_aw_valid = auto_in_aw_valid; // @[Xbar.scala 298:22]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id; // @[Xbar.scala 95:47]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_len = auto_in_aw_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_size = auto_in_aw_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_burst = auto_in_aw_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_lock = auto_in_aw_bits_lock; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_cache = auto_in_aw_bits_cache; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_prot = auto_in_aw_bits_prot; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_qos = auto_in_aw_bits_qos; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_w_valid = auto_in_w_valid; // @[Xbar.scala 242:40]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_w_bits_strb = auto_in_w_bits_strb; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_b_ready = auto_in_b_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_valid = auto_in_ar_valid; // @[Xbar.scala 298:22]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id; // @[Xbar.scala 96:47]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_len = auto_in_ar_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_burst = auto_in_ar_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_lock = auto_in_ar_bits_lock; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_cache = auto_in_ar_bits_cache; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_prot = auto_in_ar_bits_prot; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_qos = auto_in_ar_bits_qos; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_r_ready = auto_in_r_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_awOut_0_io_enq_bits_T_4 & ~(_awOut_0_io_enq_bits_T_1 | auto_in_aw_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:278 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 278:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_awOut_0_io_enq_bits_T_1 | auto_in_aw_valid) & _awOut_0_io_enq_bits_T_4) begin
          $fatal; // @[Xbar.scala 278:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_awOut_0_io_enq_bits_T_4 & ~(_T_1 | auto_in_ar_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:278 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 278:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_1 | auto_in_ar_valid) & _awOut_0_io_enq_bits_T_4) begin
          $fatal; // @[Xbar.scala 278:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_awOut_0_io_enq_bits_T_4 & ~(_T_14 | auto_out_r_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:278 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 278:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_14 | auto_out_r_valid) & _awOut_0_io_enq_bits_T_4) begin
          $fatal; // @[Xbar.scala 278:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_awOut_0_io_enq_bits_T_4 & ~(_T_26 | auto_out_b_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:278 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 278:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_26 | auto_out_b_valid) & _awOut_0_io_enq_bits_T_4) begin
          $fatal; // @[Xbar.scala 278:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_23(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [5:0]  io_enq_bits_id,
  input  [33:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_len,
  input  [2:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_burst,
  input         io_enq_bits_lock,
  input  [3:0]  io_enq_bits_cache,
  input  [2:0]  io_enq_bits_prot,
  input  [3:0]  io_enq_bits_qos,
  input         io_deq_ready,
  output        io_deq_valid,
  output [5:0]  io_deq_bits_id,
  output [33:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_len,
  output [2:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_burst,
  output        io_deq_bits_lock,
  output [3:0]  io_deq_bits_cache,
  output [2:0]  io_deq_bits_prot,
  output [3:0]  io_deq_bits_qos
);
  reg [5:0] ram_id [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [5:0] ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [5:0] ram_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [33:0] ram_addr [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_addr_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_addr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [33:0] ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [33:0] ram_addr_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_addr_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_addr_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_addr_MPORT_en; // @[Decoupled.scala 273:95]
  reg [7:0] ram_len [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_len_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_len_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [7:0] ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [7:0] ram_len_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_len_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_len_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_len_MPORT_en; // @[Decoupled.scala 273:95]
  reg [2:0] ram_size [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_size_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_burst [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_burst_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_burst_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_burst_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_burst_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_burst_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_burst_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_lock [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_lock_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_lock_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_lock_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_lock_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_lock_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_lock_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_lock_MPORT_en; // @[Decoupled.scala 273:95]
  reg [3:0] ram_cache [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_cache_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_cache_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [3:0] ram_cache_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [3:0] ram_cache_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_cache_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_cache_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_cache_MPORT_en; // @[Decoupled.scala 273:95]
  reg [2:0] ram_prot [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_prot_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_prot_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [2:0] ram_prot_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_prot_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_prot_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_prot_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_prot_MPORT_en; // @[Decoupled.scala 273:95]
  reg [3:0] ram_qos [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_qos_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_qos_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [3:0] ram_qos_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [3:0] ram_qos_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_qos_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_qos_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_qos_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = enq_ptr_value;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_addr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_addr_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = enq_ptr_value;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_len_io_deq_bits_MPORT_en = 1'h1;
  assign ram_len_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_len_io_deq_bits_MPORT_data = ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_len_MPORT_data = io_enq_bits_len;
  assign ram_len_MPORT_addr = enq_ptr_value;
  assign ram_len_MPORT_mask = 1'h1;
  assign ram_len_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = enq_ptr_value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_burst_io_deq_bits_MPORT_en = 1'h1;
  assign ram_burst_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_burst_io_deq_bits_MPORT_data = ram_burst[ram_burst_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_burst_MPORT_data = io_enq_bits_burst;
  assign ram_burst_MPORT_addr = enq_ptr_value;
  assign ram_burst_MPORT_mask = 1'h1;
  assign ram_burst_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_lock_io_deq_bits_MPORT_en = 1'h1;
  assign ram_lock_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_lock_io_deq_bits_MPORT_data = ram_lock[ram_lock_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_lock_MPORT_data = io_enq_bits_lock;
  assign ram_lock_MPORT_addr = enq_ptr_value;
  assign ram_lock_MPORT_mask = 1'h1;
  assign ram_lock_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_cache_io_deq_bits_MPORT_en = 1'h1;
  assign ram_cache_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_cache_io_deq_bits_MPORT_data = ram_cache[ram_cache_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_cache_MPORT_data = io_enq_bits_cache;
  assign ram_cache_MPORT_addr = enq_ptr_value;
  assign ram_cache_MPORT_mask = 1'h1;
  assign ram_cache_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_prot_io_deq_bits_MPORT_en = 1'h1;
  assign ram_prot_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_prot_io_deq_bits_MPORT_data = ram_prot[ram_prot_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_prot_MPORT_data = io_enq_bits_prot;
  assign ram_prot_MPORT_addr = enq_ptr_value;
  assign ram_prot_MPORT_mask = 1'h1;
  assign ram_prot_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_qos_io_deq_bits_MPORT_en = 1'h1;
  assign ram_qos_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_qos_io_deq_bits_MPORT_data = ram_qos[ram_qos_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_qos_MPORT_data = io_enq_bits_qos;
  assign ram_qos_MPORT_addr = enq_ptr_value;
  assign ram_qos_MPORT_mask = 1'h1;
  assign ram_qos_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_id = ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_addr = ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_len = ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_burst = ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_lock = ram_lock_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_cache = ram_cache_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_prot = ram_prot_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_qos = ram_qos_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_len_MPORT_en & ram_len_MPORT_mask) begin
      ram_len[ram_len_MPORT_addr] <= ram_len_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_burst_MPORT_en & ram_burst_MPORT_mask) begin
      ram_burst[ram_burst_MPORT_addr] <= ram_burst_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_lock_MPORT_en & ram_lock_MPORT_mask) begin
      ram_lock[ram_lock_MPORT_addr] <= ram_lock_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_cache_MPORT_en & ram_cache_MPORT_mask) begin
      ram_cache[ram_cache_MPORT_addr] <= ram_cache_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_prot_MPORT_en & ram_prot_MPORT_mask) begin
      ram_prot[ram_prot_MPORT_addr] <= ram_prot_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_qos_MPORT_en & ram_qos_MPORT_mask) begin
      ram_qos[ram_qos_MPORT_addr] <= ram_qos_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
endmodule
module Queue_25(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [5:0] io_enq_bits_id,
  input  [1:0] io_enq_bits_resp,
  input        io_deq_ready,
  output       io_deq_valid,
  output [5:0] io_deq_bits_id,
  output [1:0] io_deq_bits_resp
);
  reg [5:0] ram_id [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [5:0] ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [5:0] ram_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_resp [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_resp_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_resp_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_resp_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = enq_ptr_value;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_resp_io_deq_bits_MPORT_en = 1'h1;
  assign ram_resp_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_resp_io_deq_bits_MPORT_data = ram_resp[ram_resp_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_resp_MPORT_data = io_enq_bits_resp;
  assign ram_resp_MPORT_addr = enq_ptr_value;
  assign ram_resp_MPORT_mask = 1'h1;
  assign ram_resp_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_id = ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_resp = ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_resp_MPORT_en & ram_resp_MPORT_mask) begin
      ram_resp[ram_resp_MPORT_addr] <= ram_resp_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
endmodule
module Queue_27(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [5:0]   io_enq_bits_id,
  input  [511:0] io_enq_bits_data,
  input  [1:0]   io_enq_bits_resp,
  input          io_enq_bits_last,
  input          io_deq_ready,
  output         io_deq_valid,
  output [5:0]   io_deq_bits_id,
  output [511:0] io_deq_bits_data,
  output [1:0]   io_deq_bits_resp,
  output         io_deq_bits_last
);
  reg [5:0] ram_id [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [5:0] ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [5:0] ram_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [511:0] ram_data [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [511:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [511:0] ram_data_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_resp [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_resp_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_resp_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_resp_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_last [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = enq_ptr_value;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_resp_io_deq_bits_MPORT_en = 1'h1;
  assign ram_resp_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_resp_io_deq_bits_MPORT_data = ram_resp[ram_resp_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_resp_MPORT_data = io_enq_bits_resp;
  assign ram_resp_MPORT_addr = enq_ptr_value;
  assign ram_resp_MPORT_mask = 1'h1;
  assign ram_resp_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_last_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_last_io_deq_bits_MPORT_data = ram_last[ram_last_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_last_MPORT_data = io_enq_bits_last;
  assign ram_last_MPORT_addr = enq_ptr_value;
  assign ram_last_MPORT_mask = 1'h1;
  assign ram_last_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_id = ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_resp = ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_last = ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_resp_MPORT_en & ram_resp_MPORT_mask) begin
      ram_resp[ram_resp_MPORT_addr] <= ram_resp_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_last_MPORT_en & ram_last_MPORT_mask) begin
      ram_last[ram_last_MPORT_addr] <= ram_last_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
endmodule
module AXI4Buffer_2(
  input          clock,
  input          reset,
  output         auto_in_aw_ready,
  input          auto_in_aw_valid,
  input  [5:0]   auto_in_aw_bits_id,
  input  [33:0]  auto_in_aw_bits_addr,
  input  [7:0]   auto_in_aw_bits_len,
  input  [2:0]   auto_in_aw_bits_size,
  input  [1:0]   auto_in_aw_bits_burst,
  input          auto_in_aw_bits_lock,
  input  [3:0]   auto_in_aw_bits_cache,
  input  [2:0]   auto_in_aw_bits_prot,
  input  [3:0]   auto_in_aw_bits_qos,
  output         auto_in_w_ready,
  input          auto_in_w_valid,
  input  [511:0] auto_in_w_bits_data,
  input  [63:0]  auto_in_w_bits_strb,
  input          auto_in_w_bits_last,
  input          auto_in_b_ready,
  output         auto_in_b_valid,
  output [5:0]   auto_in_b_bits_id,
  output [1:0]   auto_in_b_bits_resp,
  output         auto_in_ar_ready,
  input          auto_in_ar_valid,
  input  [5:0]   auto_in_ar_bits_id,
  input  [33:0]  auto_in_ar_bits_addr,
  input  [7:0]   auto_in_ar_bits_len,
  input  [2:0]   auto_in_ar_bits_size,
  input  [1:0]   auto_in_ar_bits_burst,
  input          auto_in_ar_bits_lock,
  input  [3:0]   auto_in_ar_bits_cache,
  input  [2:0]   auto_in_ar_bits_prot,
  input  [3:0]   auto_in_ar_bits_qos,
  input          auto_in_r_ready,
  output         auto_in_r_valid,
  output [5:0]   auto_in_r_bits_id,
  output [511:0] auto_in_r_bits_data,
  output [1:0]   auto_in_r_bits_resp,
  output         auto_in_r_bits_last,
  input          auto_out_aw_ready,
  output         auto_out_aw_valid,
  output [5:0]   auto_out_aw_bits_id,
  output [33:0]  auto_out_aw_bits_addr,
  output [7:0]   auto_out_aw_bits_len,
  output [2:0]   auto_out_aw_bits_size,
  output [1:0]   auto_out_aw_bits_burst,
  output         auto_out_aw_bits_lock,
  output [3:0]   auto_out_aw_bits_cache,
  output [2:0]   auto_out_aw_bits_prot,
  output [3:0]   auto_out_aw_bits_qos,
  input          auto_out_w_ready,
  output         auto_out_w_valid,
  output [511:0] auto_out_w_bits_data,
  output [63:0]  auto_out_w_bits_strb,
  output         auto_out_w_bits_last,
  output         auto_out_b_ready,
  input          auto_out_b_valid,
  input  [5:0]   auto_out_b_bits_id,
  input  [1:0]   auto_out_b_bits_resp,
  input          auto_out_ar_ready,
  output         auto_out_ar_valid,
  output [5:0]   auto_out_ar_bits_id,
  output [33:0]  auto_out_ar_bits_addr,
  output [7:0]   auto_out_ar_bits_len,
  output [2:0]   auto_out_ar_bits_size,
  output [1:0]   auto_out_ar_bits_burst,
  output         auto_out_ar_bits_lock,
  output [3:0]   auto_out_ar_bits_cache,
  output [2:0]   auto_out_ar_bits_prot,
  output [3:0]   auto_out_ar_bits_qos,
  output         auto_out_r_ready,
  input          auto_out_r_valid,
  input  [5:0]   auto_out_r_bits_id,
  input  [511:0] auto_out_r_bits_data,
  input  [1:0]   auto_out_r_bits_resp,
  input          auto_out_r_bits_last
);
  wire  x1_aw_deq_clock; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_reset; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [5:0] x1_aw_deq_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire [33:0] x1_aw_deq_io_enq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] x1_aw_deq_io_enq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] x1_aw_deq_io_enq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] x1_aw_deq_io_enq_bits_burst; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_enq_bits_lock; // @[Decoupled.scala 375:21]
  wire [3:0] x1_aw_deq_io_enq_bits_cache; // @[Decoupled.scala 375:21]
  wire [2:0] x1_aw_deq_io_enq_bits_prot; // @[Decoupled.scala 375:21]
  wire [3:0] x1_aw_deq_io_enq_bits_qos; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [5:0] x1_aw_deq_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [33:0] x1_aw_deq_io_deq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] x1_aw_deq_io_deq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] x1_aw_deq_io_deq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] x1_aw_deq_io_deq_bits_burst; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_deq_bits_lock; // @[Decoupled.scala 375:21]
  wire [3:0] x1_aw_deq_io_deq_bits_cache; // @[Decoupled.scala 375:21]
  wire [2:0] x1_aw_deq_io_deq_bits_prot; // @[Decoupled.scala 375:21]
  wire [3:0] x1_aw_deq_io_deq_bits_qos; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_clock; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_reset; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [511:0] x1_w_deq_io_enq_bits_data; // @[Decoupled.scala 375:21]
  wire [63:0] x1_w_deq_io_enq_bits_strb; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_enq_bits_last; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [511:0] x1_w_deq_io_deq_bits_data; // @[Decoupled.scala 375:21]
  wire [63:0] x1_w_deq_io_deq_bits_strb; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_deq_bits_last; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_clock; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_reset; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [5:0] bundleIn_0_b_deq_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire [1:0] bundleIn_0_b_deq_io_enq_bits_resp; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [5:0] bundleIn_0_b_deq_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [1:0] bundleIn_0_b_deq_io_deq_bits_resp; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_clock; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_reset; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [5:0] x1_ar_deq_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire [33:0] x1_ar_deq_io_enq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] x1_ar_deq_io_enq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] x1_ar_deq_io_enq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] x1_ar_deq_io_enq_bits_burst; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_enq_bits_lock; // @[Decoupled.scala 375:21]
  wire [3:0] x1_ar_deq_io_enq_bits_cache; // @[Decoupled.scala 375:21]
  wire [2:0] x1_ar_deq_io_enq_bits_prot; // @[Decoupled.scala 375:21]
  wire [3:0] x1_ar_deq_io_enq_bits_qos; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [5:0] x1_ar_deq_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [33:0] x1_ar_deq_io_deq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] x1_ar_deq_io_deq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] x1_ar_deq_io_deq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] x1_ar_deq_io_deq_bits_burst; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_deq_bits_lock; // @[Decoupled.scala 375:21]
  wire [3:0] x1_ar_deq_io_deq_bits_cache; // @[Decoupled.scala 375:21]
  wire [2:0] x1_ar_deq_io_deq_bits_prot; // @[Decoupled.scala 375:21]
  wire [3:0] x1_ar_deq_io_deq_bits_qos; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_clock; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_reset; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [5:0] bundleIn_0_r_deq_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire [511:0] bundleIn_0_r_deq_io_enq_bits_data; // @[Decoupled.scala 375:21]
  wire [1:0] bundleIn_0_r_deq_io_enq_bits_resp; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_enq_bits_last; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [5:0] bundleIn_0_r_deq_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [511:0] bundleIn_0_r_deq_io_deq_bits_data; // @[Decoupled.scala 375:21]
  wire [1:0] bundleIn_0_r_deq_io_deq_bits_resp; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_deq_bits_last; // @[Decoupled.scala 375:21]
  Queue_23 x1_aw_deq ( // @[Decoupled.scala 375:21]
    .clock(x1_aw_deq_clock),
    .reset(x1_aw_deq_reset),
    .io_enq_ready(x1_aw_deq_io_enq_ready),
    .io_enq_valid(x1_aw_deq_io_enq_valid),
    .io_enq_bits_id(x1_aw_deq_io_enq_bits_id),
    .io_enq_bits_addr(x1_aw_deq_io_enq_bits_addr),
    .io_enq_bits_len(x1_aw_deq_io_enq_bits_len),
    .io_enq_bits_size(x1_aw_deq_io_enq_bits_size),
    .io_enq_bits_burst(x1_aw_deq_io_enq_bits_burst),
    .io_enq_bits_lock(x1_aw_deq_io_enq_bits_lock),
    .io_enq_bits_cache(x1_aw_deq_io_enq_bits_cache),
    .io_enq_bits_prot(x1_aw_deq_io_enq_bits_prot),
    .io_enq_bits_qos(x1_aw_deq_io_enq_bits_qos),
    .io_deq_ready(x1_aw_deq_io_deq_ready),
    .io_deq_valid(x1_aw_deq_io_deq_valid),
    .io_deq_bits_id(x1_aw_deq_io_deq_bits_id),
    .io_deq_bits_addr(x1_aw_deq_io_deq_bits_addr),
    .io_deq_bits_len(x1_aw_deq_io_deq_bits_len),
    .io_deq_bits_size(x1_aw_deq_io_deq_bits_size),
    .io_deq_bits_burst(x1_aw_deq_io_deq_bits_burst),
    .io_deq_bits_lock(x1_aw_deq_io_deq_bits_lock),
    .io_deq_bits_cache(x1_aw_deq_io_deq_bits_cache),
    .io_deq_bits_prot(x1_aw_deq_io_deq_bits_prot),
    .io_deq_bits_qos(x1_aw_deq_io_deq_bits_qos)
  );
  Queue_7 x1_w_deq ( // @[Decoupled.scala 375:21]
    .clock(x1_w_deq_clock),
    .reset(x1_w_deq_reset),
    .io_enq_ready(x1_w_deq_io_enq_ready),
    .io_enq_valid(x1_w_deq_io_enq_valid),
    .io_enq_bits_data(x1_w_deq_io_enq_bits_data),
    .io_enq_bits_strb(x1_w_deq_io_enq_bits_strb),
    .io_enq_bits_last(x1_w_deq_io_enq_bits_last),
    .io_deq_ready(x1_w_deq_io_deq_ready),
    .io_deq_valid(x1_w_deq_io_deq_valid),
    .io_deq_bits_data(x1_w_deq_io_deq_bits_data),
    .io_deq_bits_strb(x1_w_deq_io_deq_bits_strb),
    .io_deq_bits_last(x1_w_deq_io_deq_bits_last)
  );
  Queue_25 bundleIn_0_b_deq ( // @[Decoupled.scala 375:21]
    .clock(bundleIn_0_b_deq_clock),
    .reset(bundleIn_0_b_deq_reset),
    .io_enq_ready(bundleIn_0_b_deq_io_enq_ready),
    .io_enq_valid(bundleIn_0_b_deq_io_enq_valid),
    .io_enq_bits_id(bundleIn_0_b_deq_io_enq_bits_id),
    .io_enq_bits_resp(bundleIn_0_b_deq_io_enq_bits_resp),
    .io_deq_ready(bundleIn_0_b_deq_io_deq_ready),
    .io_deq_valid(bundleIn_0_b_deq_io_deq_valid),
    .io_deq_bits_id(bundleIn_0_b_deq_io_deq_bits_id),
    .io_deq_bits_resp(bundleIn_0_b_deq_io_deq_bits_resp)
  );
  Queue_23 x1_ar_deq ( // @[Decoupled.scala 375:21]
    .clock(x1_ar_deq_clock),
    .reset(x1_ar_deq_reset),
    .io_enq_ready(x1_ar_deq_io_enq_ready),
    .io_enq_valid(x1_ar_deq_io_enq_valid),
    .io_enq_bits_id(x1_ar_deq_io_enq_bits_id),
    .io_enq_bits_addr(x1_ar_deq_io_enq_bits_addr),
    .io_enq_bits_len(x1_ar_deq_io_enq_bits_len),
    .io_enq_bits_size(x1_ar_deq_io_enq_bits_size),
    .io_enq_bits_burst(x1_ar_deq_io_enq_bits_burst),
    .io_enq_bits_lock(x1_ar_deq_io_enq_bits_lock),
    .io_enq_bits_cache(x1_ar_deq_io_enq_bits_cache),
    .io_enq_bits_prot(x1_ar_deq_io_enq_bits_prot),
    .io_enq_bits_qos(x1_ar_deq_io_enq_bits_qos),
    .io_deq_ready(x1_ar_deq_io_deq_ready),
    .io_deq_valid(x1_ar_deq_io_deq_valid),
    .io_deq_bits_id(x1_ar_deq_io_deq_bits_id),
    .io_deq_bits_addr(x1_ar_deq_io_deq_bits_addr),
    .io_deq_bits_len(x1_ar_deq_io_deq_bits_len),
    .io_deq_bits_size(x1_ar_deq_io_deq_bits_size),
    .io_deq_bits_burst(x1_ar_deq_io_deq_bits_burst),
    .io_deq_bits_lock(x1_ar_deq_io_deq_bits_lock),
    .io_deq_bits_cache(x1_ar_deq_io_deq_bits_cache),
    .io_deq_bits_prot(x1_ar_deq_io_deq_bits_prot),
    .io_deq_bits_qos(x1_ar_deq_io_deq_bits_qos)
  );
  Queue_27 bundleIn_0_r_deq ( // @[Decoupled.scala 375:21]
    .clock(bundleIn_0_r_deq_clock),
    .reset(bundleIn_0_r_deq_reset),
    .io_enq_ready(bundleIn_0_r_deq_io_enq_ready),
    .io_enq_valid(bundleIn_0_r_deq_io_enq_valid),
    .io_enq_bits_id(bundleIn_0_r_deq_io_enq_bits_id),
    .io_enq_bits_data(bundleIn_0_r_deq_io_enq_bits_data),
    .io_enq_bits_resp(bundleIn_0_r_deq_io_enq_bits_resp),
    .io_enq_bits_last(bundleIn_0_r_deq_io_enq_bits_last),
    .io_deq_ready(bundleIn_0_r_deq_io_deq_ready),
    .io_deq_valid(bundleIn_0_r_deq_io_deq_valid),
    .io_deq_bits_id(bundleIn_0_r_deq_io_deq_bits_id),
    .io_deq_bits_data(bundleIn_0_r_deq_io_deq_bits_data),
    .io_deq_bits_resp(bundleIn_0_r_deq_io_deq_bits_resp),
    .io_deq_bits_last(bundleIn_0_r_deq_io_deq_bits_last)
  );
  assign auto_in_aw_ready = x1_aw_deq_io_enq_ready; // @[Nodes.scala 1215:84 Decoupled.scala 379:17]
  assign auto_in_w_ready = x1_w_deq_io_enq_ready; // @[Nodes.scala 1215:84 Decoupled.scala 379:17]
  assign auto_in_b_valid = bundleIn_0_b_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_in_b_bits_id = bundleIn_0_b_deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_b_bits_resp = bundleIn_0_b_deq_io_deq_bits_resp; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_ar_ready = x1_ar_deq_io_enq_ready; // @[Nodes.scala 1215:84 Decoupled.scala 379:17]
  assign auto_in_r_valid = bundleIn_0_r_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_in_r_bits_id = bundleIn_0_r_deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_r_bits_data = bundleIn_0_r_deq_io_deq_bits_data; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_r_bits_resp = bundleIn_0_r_deq_io_deq_bits_resp; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_r_bits_last = bundleIn_0_r_deq_io_deq_bits_last; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_valid = x1_aw_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_out_aw_bits_id = x1_aw_deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_addr = x1_aw_deq_io_deq_bits_addr; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_len = x1_aw_deq_io_deq_bits_len; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_size = x1_aw_deq_io_deq_bits_size; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_burst = x1_aw_deq_io_deq_bits_burst; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_lock = x1_aw_deq_io_deq_bits_lock; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_cache = x1_aw_deq_io_deq_bits_cache; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_prot = x1_aw_deq_io_deq_bits_prot; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_qos = x1_aw_deq_io_deq_bits_qos; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_w_valid = x1_w_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_out_w_bits_data = x1_w_deq_io_deq_bits_data; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_w_bits_strb = x1_w_deq_io_deq_bits_strb; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_w_bits_last = x1_w_deq_io_deq_bits_last; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_b_ready = bundleIn_0_b_deq_io_enq_ready; // @[Nodes.scala 1212:84 Decoupled.scala 379:17]
  assign auto_out_ar_valid = x1_ar_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_out_ar_bits_id = x1_ar_deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_addr = x1_ar_deq_io_deq_bits_addr; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_len = x1_ar_deq_io_deq_bits_len; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_size = x1_ar_deq_io_deq_bits_size; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_burst = x1_ar_deq_io_deq_bits_burst; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_lock = x1_ar_deq_io_deq_bits_lock; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_cache = x1_ar_deq_io_deq_bits_cache; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_prot = x1_ar_deq_io_deq_bits_prot; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_qos = x1_ar_deq_io_deq_bits_qos; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_r_ready = bundleIn_0_r_deq_io_enq_ready; // @[Nodes.scala 1212:84 Decoupled.scala 379:17]
  assign x1_aw_deq_clock = clock;
  assign x1_aw_deq_reset = reset;
  assign x1_aw_deq_io_enq_valid = auto_in_aw_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_id = auto_in_aw_bits_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_addr = auto_in_aw_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_len = auto_in_aw_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_size = auto_in_aw_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_burst = auto_in_aw_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_lock = auto_in_aw_bits_lock; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_cache = auto_in_aw_bits_cache; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_prot = auto_in_aw_bits_prot; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_qos = auto_in_aw_bits_qos; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_deq_ready = auto_out_aw_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign x1_w_deq_clock = clock;
  assign x1_w_deq_reset = reset;
  assign x1_w_deq_io_enq_valid = auto_in_w_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_w_deq_io_enq_bits_data = auto_in_w_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_w_deq_io_enq_bits_strb = auto_in_w_bits_strb; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_w_deq_io_enq_bits_last = auto_in_w_bits_last; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_w_deq_io_deq_ready = auto_out_w_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_b_deq_clock = clock;
  assign bundleIn_0_b_deq_reset = reset;
  assign bundleIn_0_b_deq_io_enq_valid = auto_out_b_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_b_deq_io_enq_bits_id = auto_out_b_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_b_deq_io_enq_bits_resp = auto_out_b_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_b_deq_io_deq_ready = auto_in_b_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_clock = clock;
  assign x1_ar_deq_reset = reset;
  assign x1_ar_deq_io_enq_valid = auto_in_ar_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_id = auto_in_ar_bits_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_addr = auto_in_ar_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_len = auto_in_ar_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_size = auto_in_ar_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_burst = auto_in_ar_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_lock = auto_in_ar_bits_lock; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_cache = auto_in_ar_bits_cache; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_prot = auto_in_ar_bits_prot; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_qos = auto_in_ar_bits_qos; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_deq_ready = auto_out_ar_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_clock = clock;
  assign bundleIn_0_r_deq_reset = reset;
  assign bundleIn_0_r_deq_io_enq_valid = auto_out_r_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_enq_bits_id = auto_out_r_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_enq_bits_data = auto_out_r_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_enq_bits_resp = auto_out_r_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_enq_bits_last = auto_out_r_bits_last; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_deq_ready = auto_in_r_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
endmodule
module Queue_33(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [6:0] io_enq_bits_tl_state_source,
  input  [1:0] io_enq_bits_extra_id,
  input        io_deq_ready,
  output       io_deq_valid,
  output [6:0] io_deq_bits_tl_state_source,
  output [1:0] io_deq_bits_extra_id
);
  reg [6:0] ram_tl_state_source [0:3]; // @[Decoupled.scala 273:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_tl_state_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [6:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [6:0] ram_tl_state_source_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_tl_state_source_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tl_state_source_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_tl_state_source_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_extra_id [0:3]; // @[Decoupled.scala 273:95]
  wire  ram_extra_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_extra_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_extra_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_extra_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_extra_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_extra_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = enq_ptr_value;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_extra_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_extra_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_extra_id_io_deq_bits_MPORT_data = ram_extra_id[ram_extra_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_extra_id_MPORT_data = io_enq_bits_extra_id;
  assign ram_extra_id_MPORT_addr = enq_ptr_value;
  assign ram_extra_id_MPORT_mask = 1'h1;
  assign ram_extra_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_extra_id = ram_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_extra_id_MPORT_en & ram_extra_id_MPORT_mask) begin
      ram_extra_id[ram_extra_id_MPORT_addr] <= ram_extra_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
endmodule
module Queue_35(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [6:0] io_enq_bits_tl_state_source,
  input  [1:0] io_enq_bits_extra_id,
  input        io_deq_ready,
  output       io_deq_valid,
  output [6:0] io_deq_bits_tl_state_source,
  output [1:0] io_deq_bits_extra_id
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_GARBAGE_ASSIGN
  reg [6:0] ram_tl_state_source [0:2]; // @[Decoupled.scala 273:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_tl_state_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [6:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [6:0] ram_tl_state_source_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_tl_state_source_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tl_state_source_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_tl_state_source_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_extra_id [0:2]; // @[Decoupled.scala 273:95]
  wire  ram_extra_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_extra_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_extra_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_extra_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_extra_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_extra_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire  wrap = enq_ptr_value == 2'h2; // @[Counter.scala 73:24]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire  wrap_1 = deq_ptr_value == 2'h2; // @[Counter.scala 73:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `else
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_0[6:0]
     : ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = enq_ptr_value;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_extra_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_extra_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_extra_id_io_deq_bits_MPORT_data = ram_extra_id[ram_extra_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `else
  assign ram_extra_id_io_deq_bits_MPORT_data = ram_extra_id_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_1[1:0] :
    ram_extra_id[ram_extra_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_extra_id_MPORT_data = io_enq_bits_extra_id;
  assign ram_extra_id_MPORT_addr = enq_ptr_value;
  assign ram_extra_id_MPORT_mask = 1'h1;
  assign ram_extra_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_extra_id = ram_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_extra_id_MPORT_en & ram_extra_id_MPORT_mask) begin
      ram_extra_id[ram_extra_id_MPORT_addr] <= ram_extra_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      if (wrap) begin // @[Counter.scala 87:20]
        enq_ptr_value <= 2'h0; // @[Counter.scala 87:28]
      end else begin
        enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
      end
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      if (wrap_1) begin // @[Counter.scala 87:20]
        deq_ptr_value <= 2'h0; // @[Counter.scala 87:28]
      end else begin
        deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
      end
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_0 = {1{`RANDOM}};
  _RAND_1 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4UserYanker(
  input          clock,
  input          reset,
  output         auto_in_aw_ready,
  input          auto_in_aw_valid,
  input  [5:0]   auto_in_aw_bits_id,
  input  [33:0]  auto_in_aw_bits_addr,
  input  [7:0]   auto_in_aw_bits_len,
  input  [2:0]   auto_in_aw_bits_size,
  input  [1:0]   auto_in_aw_bits_burst,
  input          auto_in_aw_bits_lock,
  input  [3:0]   auto_in_aw_bits_cache,
  input  [2:0]   auto_in_aw_bits_prot,
  input  [3:0]   auto_in_aw_bits_qos,
  input  [6:0]   auto_in_aw_bits_echo_tl_state_source,
  input  [1:0]   auto_in_aw_bits_echo_extra_id,
  output         auto_in_w_ready,
  input          auto_in_w_valid,
  input  [511:0] auto_in_w_bits_data,
  input  [63:0]  auto_in_w_bits_strb,
  input          auto_in_w_bits_last,
  input          auto_in_b_ready,
  output         auto_in_b_valid,
  output [5:0]   auto_in_b_bits_id,
  output [1:0]   auto_in_b_bits_resp,
  output [6:0]   auto_in_b_bits_echo_tl_state_source,
  output [1:0]   auto_in_b_bits_echo_extra_id,
  output         auto_in_ar_ready,
  input          auto_in_ar_valid,
  input  [5:0]   auto_in_ar_bits_id,
  input  [33:0]  auto_in_ar_bits_addr,
  input  [7:0]   auto_in_ar_bits_len,
  input  [2:0]   auto_in_ar_bits_size,
  input  [1:0]   auto_in_ar_bits_burst,
  input          auto_in_ar_bits_lock,
  input  [3:0]   auto_in_ar_bits_cache,
  input  [2:0]   auto_in_ar_bits_prot,
  input  [3:0]   auto_in_ar_bits_qos,
  input  [6:0]   auto_in_ar_bits_echo_tl_state_source,
  input  [1:0]   auto_in_ar_bits_echo_extra_id,
  input          auto_in_r_ready,
  output         auto_in_r_valid,
  output [5:0]   auto_in_r_bits_id,
  output [511:0] auto_in_r_bits_data,
  output [1:0]   auto_in_r_bits_resp,
  output [6:0]   auto_in_r_bits_echo_tl_state_source,
  output [1:0]   auto_in_r_bits_echo_extra_id,
  output         auto_in_r_bits_last,
  input          auto_out_aw_ready,
  output         auto_out_aw_valid,
  output [5:0]   auto_out_aw_bits_id,
  output [33:0]  auto_out_aw_bits_addr,
  output [7:0]   auto_out_aw_bits_len,
  output [2:0]   auto_out_aw_bits_size,
  output [1:0]   auto_out_aw_bits_burst,
  output         auto_out_aw_bits_lock,
  output [3:0]   auto_out_aw_bits_cache,
  output [2:0]   auto_out_aw_bits_prot,
  output [3:0]   auto_out_aw_bits_qos,
  input          auto_out_w_ready,
  output         auto_out_w_valid,
  output [511:0] auto_out_w_bits_data,
  output [63:0]  auto_out_w_bits_strb,
  output         auto_out_w_bits_last,
  output         auto_out_b_ready,
  input          auto_out_b_valid,
  input  [5:0]   auto_out_b_bits_id,
  input  [1:0]   auto_out_b_bits_resp,
  input          auto_out_ar_ready,
  output         auto_out_ar_valid,
  output [5:0]   auto_out_ar_bits_id,
  output [33:0]  auto_out_ar_bits_addr,
  output [7:0]   auto_out_ar_bits_len,
  output [2:0]   auto_out_ar_bits_size,
  output [1:0]   auto_out_ar_bits_burst,
  output         auto_out_ar_bits_lock,
  output [3:0]   auto_out_ar_bits_cache,
  output [2:0]   auto_out_ar_bits_prot,
  output [3:0]   auto_out_ar_bits_qos,
  output         auto_out_r_ready,
  input          auto_out_r_valid,
  input  [5:0]   auto_out_r_bits_id,
  input  [511:0] auto_out_r_bits_data,
  input  [1:0]   auto_out_r_bits_resp,
  input          auto_out_r_bits_last
);
  wire  Queue_clock; // @[UserYanker.scala 50:17]
  wire  Queue_reset; // @[UserYanker.scala 50:17]
  wire  Queue_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_1_clock; // @[UserYanker.scala 50:17]
  wire  Queue_1_reset; // @[UserYanker.scala 50:17]
  wire  Queue_1_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_1_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_1_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_1_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_1_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_1_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_1_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_1_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_2_clock; // @[UserYanker.scala 50:17]
  wire  Queue_2_reset; // @[UserYanker.scala 50:17]
  wire  Queue_2_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_2_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_2_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_2_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_2_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_2_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_2_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_2_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_3_clock; // @[UserYanker.scala 50:17]
  wire  Queue_3_reset; // @[UserYanker.scala 50:17]
  wire  Queue_3_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_3_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_3_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_3_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_3_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_3_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_3_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_3_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_4_clock; // @[UserYanker.scala 50:17]
  wire  Queue_4_reset; // @[UserYanker.scala 50:17]
  wire  Queue_4_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_4_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_4_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_4_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_4_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_4_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_4_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_4_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_5_clock; // @[UserYanker.scala 50:17]
  wire  Queue_5_reset; // @[UserYanker.scala 50:17]
  wire  Queue_5_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_5_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_5_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_5_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_5_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_5_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_5_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_5_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_6_clock; // @[UserYanker.scala 50:17]
  wire  Queue_6_reset; // @[UserYanker.scala 50:17]
  wire  Queue_6_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_6_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_6_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_6_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_6_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_6_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_6_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_6_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_7_clock; // @[UserYanker.scala 50:17]
  wire  Queue_7_reset; // @[UserYanker.scala 50:17]
  wire  Queue_7_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_7_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_7_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_7_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_7_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_7_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_7_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_7_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_8_clock; // @[UserYanker.scala 50:17]
  wire  Queue_8_reset; // @[UserYanker.scala 50:17]
  wire  Queue_8_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_8_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_8_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_8_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_8_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_8_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_8_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_8_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_9_clock; // @[UserYanker.scala 50:17]
  wire  Queue_9_reset; // @[UserYanker.scala 50:17]
  wire  Queue_9_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_9_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_9_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_9_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_9_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_9_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_9_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_9_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_10_clock; // @[UserYanker.scala 50:17]
  wire  Queue_10_reset; // @[UserYanker.scala 50:17]
  wire  Queue_10_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_10_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_10_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_10_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_10_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_10_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_10_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_10_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_11_clock; // @[UserYanker.scala 50:17]
  wire  Queue_11_reset; // @[UserYanker.scala 50:17]
  wire  Queue_11_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_11_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_11_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_11_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_11_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_11_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_11_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_11_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_12_clock; // @[UserYanker.scala 50:17]
  wire  Queue_12_reset; // @[UserYanker.scala 50:17]
  wire  Queue_12_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_12_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_12_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_12_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_12_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_12_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_12_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_12_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_13_clock; // @[UserYanker.scala 50:17]
  wire  Queue_13_reset; // @[UserYanker.scala 50:17]
  wire  Queue_13_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_13_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_13_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_13_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_13_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_13_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_13_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_13_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_14_clock; // @[UserYanker.scala 50:17]
  wire  Queue_14_reset; // @[UserYanker.scala 50:17]
  wire  Queue_14_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_14_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_14_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_14_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_14_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_14_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_14_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_14_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_15_clock; // @[UserYanker.scala 50:17]
  wire  Queue_15_reset; // @[UserYanker.scala 50:17]
  wire  Queue_15_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_15_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_15_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_15_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_15_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_15_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_15_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_15_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_16_clock; // @[UserYanker.scala 50:17]
  wire  Queue_16_reset; // @[UserYanker.scala 50:17]
  wire  Queue_16_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_16_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_16_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_16_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_16_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_16_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_16_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_16_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_17_clock; // @[UserYanker.scala 50:17]
  wire  Queue_17_reset; // @[UserYanker.scala 50:17]
  wire  Queue_17_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_17_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_17_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_17_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_17_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_17_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_17_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_17_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_18_clock; // @[UserYanker.scala 50:17]
  wire  Queue_18_reset; // @[UserYanker.scala 50:17]
  wire  Queue_18_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_18_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_18_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_18_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_18_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_18_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_18_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_18_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_19_clock; // @[UserYanker.scala 50:17]
  wire  Queue_19_reset; // @[UserYanker.scala 50:17]
  wire  Queue_19_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_19_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_19_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_19_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_19_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_19_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_19_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_19_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_20_clock; // @[UserYanker.scala 50:17]
  wire  Queue_20_reset; // @[UserYanker.scala 50:17]
  wire  Queue_20_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_20_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_20_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_20_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_20_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_20_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_20_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_20_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_21_clock; // @[UserYanker.scala 50:17]
  wire  Queue_21_reset; // @[UserYanker.scala 50:17]
  wire  Queue_21_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_21_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_21_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_21_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_21_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_21_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_21_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_21_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_22_clock; // @[UserYanker.scala 50:17]
  wire  Queue_22_reset; // @[UserYanker.scala 50:17]
  wire  Queue_22_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_22_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_22_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_22_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_22_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_22_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_22_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_22_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_23_clock; // @[UserYanker.scala 50:17]
  wire  Queue_23_reset; // @[UserYanker.scala 50:17]
  wire  Queue_23_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_23_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_23_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_23_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_23_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_23_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_23_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_23_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_24_clock; // @[UserYanker.scala 50:17]
  wire  Queue_24_reset; // @[UserYanker.scala 50:17]
  wire  Queue_24_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_24_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_24_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_24_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_24_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_24_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_24_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_24_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_25_clock; // @[UserYanker.scala 50:17]
  wire  Queue_25_reset; // @[UserYanker.scala 50:17]
  wire  Queue_25_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_25_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_25_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_25_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_25_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_25_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_25_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_25_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_26_clock; // @[UserYanker.scala 50:17]
  wire  Queue_26_reset; // @[UserYanker.scala 50:17]
  wire  Queue_26_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_26_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_26_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_26_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_26_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_26_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_26_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_26_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_27_clock; // @[UserYanker.scala 50:17]
  wire  Queue_27_reset; // @[UserYanker.scala 50:17]
  wire  Queue_27_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_27_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_27_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_27_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_27_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_27_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_27_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_27_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_28_clock; // @[UserYanker.scala 50:17]
  wire  Queue_28_reset; // @[UserYanker.scala 50:17]
  wire  Queue_28_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_28_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_28_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_28_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_28_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_28_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_28_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_28_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_29_clock; // @[UserYanker.scala 50:17]
  wire  Queue_29_reset; // @[UserYanker.scala 50:17]
  wire  Queue_29_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_29_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_29_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_29_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_29_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_29_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_29_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_29_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_30_clock; // @[UserYanker.scala 50:17]
  wire  Queue_30_reset; // @[UserYanker.scala 50:17]
  wire  Queue_30_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_30_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_30_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_30_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_30_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_30_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_30_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_30_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_31_clock; // @[UserYanker.scala 50:17]
  wire  Queue_31_reset; // @[UserYanker.scala 50:17]
  wire  Queue_31_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_31_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_31_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_31_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_31_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_31_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_31_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_31_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_32_clock; // @[UserYanker.scala 50:17]
  wire  Queue_32_reset; // @[UserYanker.scala 50:17]
  wire  Queue_32_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_32_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_32_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_32_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_32_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_32_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_32_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_32_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_33_clock; // @[UserYanker.scala 50:17]
  wire  Queue_33_reset; // @[UserYanker.scala 50:17]
  wire  Queue_33_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_33_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_33_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_33_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_33_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_33_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_33_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_33_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_34_clock; // @[UserYanker.scala 50:17]
  wire  Queue_34_reset; // @[UserYanker.scala 50:17]
  wire  Queue_34_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_34_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_34_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_34_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_34_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_34_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_34_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_34_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_35_clock; // @[UserYanker.scala 50:17]
  wire  Queue_35_reset; // @[UserYanker.scala 50:17]
  wire  Queue_35_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_35_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_35_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_35_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_35_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_35_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_35_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_35_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_36_clock; // @[UserYanker.scala 50:17]
  wire  Queue_36_reset; // @[UserYanker.scala 50:17]
  wire  Queue_36_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_36_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_36_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_36_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_36_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_36_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_36_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_36_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_37_clock; // @[UserYanker.scala 50:17]
  wire  Queue_37_reset; // @[UserYanker.scala 50:17]
  wire  Queue_37_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_37_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_37_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_37_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_37_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_37_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_37_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_37_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_38_clock; // @[UserYanker.scala 50:17]
  wire  Queue_38_reset; // @[UserYanker.scala 50:17]
  wire  Queue_38_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_38_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_38_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_38_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_38_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_38_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_38_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_38_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_39_clock; // @[UserYanker.scala 50:17]
  wire  Queue_39_reset; // @[UserYanker.scala 50:17]
  wire  Queue_39_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_39_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_39_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_39_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_39_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_39_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_39_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_39_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_40_clock; // @[UserYanker.scala 50:17]
  wire  Queue_40_reset; // @[UserYanker.scala 50:17]
  wire  Queue_40_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_40_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_40_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_40_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_40_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_40_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_40_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_40_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_41_clock; // @[UserYanker.scala 50:17]
  wire  Queue_41_reset; // @[UserYanker.scala 50:17]
  wire  Queue_41_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_41_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_41_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_41_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_41_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_41_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_41_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_41_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_42_clock; // @[UserYanker.scala 50:17]
  wire  Queue_42_reset; // @[UserYanker.scala 50:17]
  wire  Queue_42_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_42_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_42_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_42_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_42_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_42_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_42_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_42_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_43_clock; // @[UserYanker.scala 50:17]
  wire  Queue_43_reset; // @[UserYanker.scala 50:17]
  wire  Queue_43_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_43_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_43_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_43_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_43_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_43_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_43_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_43_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_44_clock; // @[UserYanker.scala 50:17]
  wire  Queue_44_reset; // @[UserYanker.scala 50:17]
  wire  Queue_44_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_44_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_44_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_44_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_44_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_44_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_44_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_44_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_45_clock; // @[UserYanker.scala 50:17]
  wire  Queue_45_reset; // @[UserYanker.scala 50:17]
  wire  Queue_45_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_45_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_45_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_45_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_45_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_45_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_45_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_45_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_46_clock; // @[UserYanker.scala 50:17]
  wire  Queue_46_reset; // @[UserYanker.scala 50:17]
  wire  Queue_46_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_46_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_46_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_46_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_46_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_46_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_46_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_46_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_47_clock; // @[UserYanker.scala 50:17]
  wire  Queue_47_reset; // @[UserYanker.scala 50:17]
  wire  Queue_47_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_47_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_47_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_47_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_47_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_47_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_47_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_47_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_48_clock; // @[UserYanker.scala 50:17]
  wire  Queue_48_reset; // @[UserYanker.scala 50:17]
  wire  Queue_48_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_48_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_48_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_48_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_48_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_48_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_48_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_48_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_49_clock; // @[UserYanker.scala 50:17]
  wire  Queue_49_reset; // @[UserYanker.scala 50:17]
  wire  Queue_49_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_49_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_49_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_49_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_49_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_49_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_49_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_49_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_50_clock; // @[UserYanker.scala 50:17]
  wire  Queue_50_reset; // @[UserYanker.scala 50:17]
  wire  Queue_50_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_50_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_50_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_50_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_50_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_50_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_50_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_50_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_51_clock; // @[UserYanker.scala 50:17]
  wire  Queue_51_reset; // @[UserYanker.scala 50:17]
  wire  Queue_51_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_51_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_51_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_51_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_51_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_51_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_51_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_51_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_52_clock; // @[UserYanker.scala 50:17]
  wire  Queue_52_reset; // @[UserYanker.scala 50:17]
  wire  Queue_52_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_52_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_52_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_52_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_52_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_52_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_52_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_52_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_53_clock; // @[UserYanker.scala 50:17]
  wire  Queue_53_reset; // @[UserYanker.scala 50:17]
  wire  Queue_53_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_53_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_53_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_53_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_53_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_53_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_53_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_53_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_54_clock; // @[UserYanker.scala 50:17]
  wire  Queue_54_reset; // @[UserYanker.scala 50:17]
  wire  Queue_54_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_54_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_54_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_54_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_54_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_54_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_54_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_54_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_55_clock; // @[UserYanker.scala 50:17]
  wire  Queue_55_reset; // @[UserYanker.scala 50:17]
  wire  Queue_55_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_55_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_55_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_55_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_55_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_55_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_55_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_55_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_56_clock; // @[UserYanker.scala 50:17]
  wire  Queue_56_reset; // @[UserYanker.scala 50:17]
  wire  Queue_56_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_56_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_56_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_56_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_56_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_56_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_56_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_56_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_57_clock; // @[UserYanker.scala 50:17]
  wire  Queue_57_reset; // @[UserYanker.scala 50:17]
  wire  Queue_57_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_57_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_57_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_57_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_57_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_57_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_57_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_57_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_58_clock; // @[UserYanker.scala 50:17]
  wire  Queue_58_reset; // @[UserYanker.scala 50:17]
  wire  Queue_58_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_58_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_58_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_58_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_58_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_58_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_58_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_58_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_59_clock; // @[UserYanker.scala 50:17]
  wire  Queue_59_reset; // @[UserYanker.scala 50:17]
  wire  Queue_59_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_59_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_59_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_59_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_59_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_59_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_59_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_59_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_60_clock; // @[UserYanker.scala 50:17]
  wire  Queue_60_reset; // @[UserYanker.scala 50:17]
  wire  Queue_60_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_60_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_60_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_60_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_60_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_60_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_60_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_60_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_61_clock; // @[UserYanker.scala 50:17]
  wire  Queue_61_reset; // @[UserYanker.scala 50:17]
  wire  Queue_61_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_61_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_61_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_61_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_61_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_61_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_61_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_61_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_62_clock; // @[UserYanker.scala 50:17]
  wire  Queue_62_reset; // @[UserYanker.scala 50:17]
  wire  Queue_62_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_62_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_62_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_62_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_62_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_62_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_62_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_62_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_63_clock; // @[UserYanker.scala 50:17]
  wire  Queue_63_reset; // @[UserYanker.scala 50:17]
  wire  Queue_63_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_63_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_63_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_63_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_63_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_63_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_63_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_63_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_64_clock; // @[UserYanker.scala 50:17]
  wire  Queue_64_reset; // @[UserYanker.scala 50:17]
  wire  Queue_64_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_64_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_64_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_64_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_64_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_64_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_64_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_64_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_65_clock; // @[UserYanker.scala 50:17]
  wire  Queue_65_reset; // @[UserYanker.scala 50:17]
  wire  Queue_65_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_65_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_65_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_65_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_65_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_65_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_65_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_65_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_66_clock; // @[UserYanker.scala 50:17]
  wire  Queue_66_reset; // @[UserYanker.scala 50:17]
  wire  Queue_66_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_66_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_66_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_66_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_66_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_66_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_66_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_66_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_67_clock; // @[UserYanker.scala 50:17]
  wire  Queue_67_reset; // @[UserYanker.scala 50:17]
  wire  Queue_67_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_67_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_67_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_67_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_67_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_67_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_67_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_67_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_68_clock; // @[UserYanker.scala 50:17]
  wire  Queue_68_reset; // @[UserYanker.scala 50:17]
  wire  Queue_68_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_68_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_68_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_68_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_68_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_68_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_68_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_68_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_69_clock; // @[UserYanker.scala 50:17]
  wire  Queue_69_reset; // @[UserYanker.scala 50:17]
  wire  Queue_69_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_69_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_69_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_69_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_69_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_69_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_69_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_69_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_70_clock; // @[UserYanker.scala 50:17]
  wire  Queue_70_reset; // @[UserYanker.scala 50:17]
  wire  Queue_70_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_70_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_70_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_70_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_70_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_70_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_70_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_70_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_71_clock; // @[UserYanker.scala 50:17]
  wire  Queue_71_reset; // @[UserYanker.scala 50:17]
  wire  Queue_71_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_71_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_71_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_71_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_71_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_71_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_71_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_71_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_72_clock; // @[UserYanker.scala 50:17]
  wire  Queue_72_reset; // @[UserYanker.scala 50:17]
  wire  Queue_72_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_72_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_72_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_72_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_72_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_72_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_72_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_72_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_73_clock; // @[UserYanker.scala 50:17]
  wire  Queue_73_reset; // @[UserYanker.scala 50:17]
  wire  Queue_73_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_73_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_73_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_73_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_73_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_73_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_73_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_73_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_74_clock; // @[UserYanker.scala 50:17]
  wire  Queue_74_reset; // @[UserYanker.scala 50:17]
  wire  Queue_74_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_74_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_74_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_74_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_74_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_74_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_74_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_74_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_75_clock; // @[UserYanker.scala 50:17]
  wire  Queue_75_reset; // @[UserYanker.scala 50:17]
  wire  Queue_75_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_75_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_75_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_75_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_75_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_75_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_75_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_75_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_76_clock; // @[UserYanker.scala 50:17]
  wire  Queue_76_reset; // @[UserYanker.scala 50:17]
  wire  Queue_76_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_76_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_76_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_76_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_76_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_76_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_76_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_76_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_77_clock; // @[UserYanker.scala 50:17]
  wire  Queue_77_reset; // @[UserYanker.scala 50:17]
  wire  Queue_77_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_77_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_77_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_77_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_77_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_77_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_77_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_77_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_78_clock; // @[UserYanker.scala 50:17]
  wire  Queue_78_reset; // @[UserYanker.scala 50:17]
  wire  Queue_78_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_78_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_78_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_78_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_78_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_78_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_78_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_78_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_79_clock; // @[UserYanker.scala 50:17]
  wire  Queue_79_reset; // @[UserYanker.scala 50:17]
  wire  Queue_79_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_79_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_79_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_79_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_79_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_79_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_79_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_79_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_80_clock; // @[UserYanker.scala 50:17]
  wire  Queue_80_reset; // @[UserYanker.scala 50:17]
  wire  Queue_80_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_80_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_80_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_80_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_80_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_80_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_80_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_80_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_81_clock; // @[UserYanker.scala 50:17]
  wire  Queue_81_reset; // @[UserYanker.scala 50:17]
  wire  Queue_81_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_81_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_81_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_81_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_81_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_81_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_81_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_81_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_82_clock; // @[UserYanker.scala 50:17]
  wire  Queue_82_reset; // @[UserYanker.scala 50:17]
  wire  Queue_82_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_82_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_82_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_82_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_82_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_82_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_82_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_82_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_83_clock; // @[UserYanker.scala 50:17]
  wire  Queue_83_reset; // @[UserYanker.scala 50:17]
  wire  Queue_83_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_83_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_83_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_83_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_83_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_83_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_83_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_83_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_84_clock; // @[UserYanker.scala 50:17]
  wire  Queue_84_reset; // @[UserYanker.scala 50:17]
  wire  Queue_84_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_84_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_84_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_84_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_84_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_84_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_84_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_84_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_85_clock; // @[UserYanker.scala 50:17]
  wire  Queue_85_reset; // @[UserYanker.scala 50:17]
  wire  Queue_85_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_85_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_85_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_85_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_85_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_85_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_85_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_85_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_86_clock; // @[UserYanker.scala 50:17]
  wire  Queue_86_reset; // @[UserYanker.scala 50:17]
  wire  Queue_86_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_86_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_86_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_86_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_86_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_86_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_86_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_86_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_87_clock; // @[UserYanker.scala 50:17]
  wire  Queue_87_reset; // @[UserYanker.scala 50:17]
  wire  Queue_87_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_87_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_87_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_87_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_87_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_87_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_87_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_87_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_88_clock; // @[UserYanker.scala 50:17]
  wire  Queue_88_reset; // @[UserYanker.scala 50:17]
  wire  Queue_88_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_88_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_88_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_88_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_88_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_88_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_88_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_88_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_89_clock; // @[UserYanker.scala 50:17]
  wire  Queue_89_reset; // @[UserYanker.scala 50:17]
  wire  Queue_89_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_89_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_89_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_89_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_89_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_89_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_89_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_89_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_90_clock; // @[UserYanker.scala 50:17]
  wire  Queue_90_reset; // @[UserYanker.scala 50:17]
  wire  Queue_90_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_90_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_90_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_90_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_90_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_90_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_90_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_90_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_91_clock; // @[UserYanker.scala 50:17]
  wire  Queue_91_reset; // @[UserYanker.scala 50:17]
  wire  Queue_91_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_91_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_91_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_91_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_91_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_91_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_91_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_91_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_92_clock; // @[UserYanker.scala 50:17]
  wire  Queue_92_reset; // @[UserYanker.scala 50:17]
  wire  Queue_92_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_92_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_92_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_92_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_92_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_92_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_92_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_92_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_93_clock; // @[UserYanker.scala 50:17]
  wire  Queue_93_reset; // @[UserYanker.scala 50:17]
  wire  Queue_93_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_93_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_93_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_93_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_93_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_93_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_93_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_93_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_94_clock; // @[UserYanker.scala 50:17]
  wire  Queue_94_reset; // @[UserYanker.scala 50:17]
  wire  Queue_94_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_94_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_94_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_94_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_94_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_94_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_94_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_94_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_95_clock; // @[UserYanker.scala 50:17]
  wire  Queue_95_reset; // @[UserYanker.scala 50:17]
  wire  Queue_95_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_95_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_95_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_95_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_95_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_95_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_95_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_95_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_96_clock; // @[UserYanker.scala 50:17]
  wire  Queue_96_reset; // @[UserYanker.scala 50:17]
  wire  Queue_96_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_96_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_96_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_96_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_96_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_96_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_96_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_96_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_97_clock; // @[UserYanker.scala 50:17]
  wire  Queue_97_reset; // @[UserYanker.scala 50:17]
  wire  Queue_97_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_97_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_97_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_97_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_97_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_97_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_97_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_97_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_98_clock; // @[UserYanker.scala 50:17]
  wire  Queue_98_reset; // @[UserYanker.scala 50:17]
  wire  Queue_98_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_98_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_98_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_98_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_98_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_98_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_98_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_98_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_99_clock; // @[UserYanker.scala 50:17]
  wire  Queue_99_reset; // @[UserYanker.scala 50:17]
  wire  Queue_99_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_99_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_99_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_99_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_99_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_99_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_99_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_99_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_100_clock; // @[UserYanker.scala 50:17]
  wire  Queue_100_reset; // @[UserYanker.scala 50:17]
  wire  Queue_100_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_100_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_100_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_100_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_100_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_100_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_100_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_100_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_101_clock; // @[UserYanker.scala 50:17]
  wire  Queue_101_reset; // @[UserYanker.scala 50:17]
  wire  Queue_101_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_101_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_101_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_101_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_101_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_101_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_101_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_101_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_102_clock; // @[UserYanker.scala 50:17]
  wire  Queue_102_reset; // @[UserYanker.scala 50:17]
  wire  Queue_102_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_102_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_102_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_102_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_102_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_102_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_102_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_102_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_103_clock; // @[UserYanker.scala 50:17]
  wire  Queue_103_reset; // @[UserYanker.scala 50:17]
  wire  Queue_103_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_103_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_103_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_103_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_103_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_103_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_103_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_103_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_104_clock; // @[UserYanker.scala 50:17]
  wire  Queue_104_reset; // @[UserYanker.scala 50:17]
  wire  Queue_104_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_104_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_104_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_104_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_104_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_104_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_104_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_104_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_105_clock; // @[UserYanker.scala 50:17]
  wire  Queue_105_reset; // @[UserYanker.scala 50:17]
  wire  Queue_105_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_105_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_105_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_105_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_105_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_105_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_105_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_105_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_106_clock; // @[UserYanker.scala 50:17]
  wire  Queue_106_reset; // @[UserYanker.scala 50:17]
  wire  Queue_106_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_106_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_106_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_106_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_106_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_106_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_106_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_106_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_107_clock; // @[UserYanker.scala 50:17]
  wire  Queue_107_reset; // @[UserYanker.scala 50:17]
  wire  Queue_107_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_107_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_107_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_107_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_107_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_107_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_107_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_107_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_108_clock; // @[UserYanker.scala 50:17]
  wire  Queue_108_reset; // @[UserYanker.scala 50:17]
  wire  Queue_108_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_108_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_108_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_108_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_108_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_108_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_108_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_108_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_109_clock; // @[UserYanker.scala 50:17]
  wire  Queue_109_reset; // @[UserYanker.scala 50:17]
  wire  Queue_109_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_109_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_109_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_109_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_109_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_109_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_109_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_109_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_110_clock; // @[UserYanker.scala 50:17]
  wire  Queue_110_reset; // @[UserYanker.scala 50:17]
  wire  Queue_110_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_110_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_110_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_110_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_110_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_110_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_110_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_110_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_111_clock; // @[UserYanker.scala 50:17]
  wire  Queue_111_reset; // @[UserYanker.scala 50:17]
  wire  Queue_111_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_111_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_111_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_111_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_111_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_111_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_111_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_111_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_112_clock; // @[UserYanker.scala 50:17]
  wire  Queue_112_reset; // @[UserYanker.scala 50:17]
  wire  Queue_112_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_112_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_112_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_112_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_112_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_112_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_112_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_112_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_113_clock; // @[UserYanker.scala 50:17]
  wire  Queue_113_reset; // @[UserYanker.scala 50:17]
  wire  Queue_113_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_113_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_113_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_113_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_113_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_113_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_113_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_113_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_114_clock; // @[UserYanker.scala 50:17]
  wire  Queue_114_reset; // @[UserYanker.scala 50:17]
  wire  Queue_114_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_114_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_114_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_114_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_114_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_114_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_114_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_114_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_115_clock; // @[UserYanker.scala 50:17]
  wire  Queue_115_reset; // @[UserYanker.scala 50:17]
  wire  Queue_115_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_115_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_115_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_115_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_115_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_115_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_115_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_115_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_116_clock; // @[UserYanker.scala 50:17]
  wire  Queue_116_reset; // @[UserYanker.scala 50:17]
  wire  Queue_116_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_116_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_116_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_116_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_116_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_116_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_116_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_116_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_117_clock; // @[UserYanker.scala 50:17]
  wire  Queue_117_reset; // @[UserYanker.scala 50:17]
  wire  Queue_117_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_117_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_117_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_117_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_117_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_117_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_117_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_117_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_118_clock; // @[UserYanker.scala 50:17]
  wire  Queue_118_reset; // @[UserYanker.scala 50:17]
  wire  Queue_118_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_118_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_118_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_118_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_118_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_118_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_118_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_118_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_119_clock; // @[UserYanker.scala 50:17]
  wire  Queue_119_reset; // @[UserYanker.scala 50:17]
  wire  Queue_119_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_119_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_119_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_119_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_119_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_119_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_119_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_119_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_120_clock; // @[UserYanker.scala 50:17]
  wire  Queue_120_reset; // @[UserYanker.scala 50:17]
  wire  Queue_120_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_120_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_120_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_120_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_120_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_120_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_120_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_120_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_121_clock; // @[UserYanker.scala 50:17]
  wire  Queue_121_reset; // @[UserYanker.scala 50:17]
  wire  Queue_121_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_121_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_121_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_121_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_121_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_121_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_121_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_121_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_122_clock; // @[UserYanker.scala 50:17]
  wire  Queue_122_reset; // @[UserYanker.scala 50:17]
  wire  Queue_122_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_122_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_122_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_122_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_122_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_122_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_122_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_122_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_123_clock; // @[UserYanker.scala 50:17]
  wire  Queue_123_reset; // @[UserYanker.scala 50:17]
  wire  Queue_123_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_123_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_123_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_123_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_123_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_123_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_123_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_123_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_124_clock; // @[UserYanker.scala 50:17]
  wire  Queue_124_reset; // @[UserYanker.scala 50:17]
  wire  Queue_124_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_124_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_124_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_124_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_124_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_124_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_124_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_124_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_125_clock; // @[UserYanker.scala 50:17]
  wire  Queue_125_reset; // @[UserYanker.scala 50:17]
  wire  Queue_125_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_125_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_125_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_125_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_125_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_125_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_125_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_125_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_126_clock; // @[UserYanker.scala 50:17]
  wire  Queue_126_reset; // @[UserYanker.scala 50:17]
  wire  Queue_126_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_126_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_126_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_126_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_126_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_126_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_126_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_126_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_127_clock; // @[UserYanker.scala 50:17]
  wire  Queue_127_reset; // @[UserYanker.scala 50:17]
  wire  Queue_127_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_127_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_127_io_enq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_127_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_127_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_127_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [6:0] Queue_127_io_deq_bits_tl_state_source; // @[UserYanker.scala 50:17]
  wire [1:0] Queue_127_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  _ar_ready_WIRE_0 = Queue_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _ar_ready_WIRE_1 = Queue_1_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_1 = 6'h1 == auto_in_ar_bits_id ? _ar_ready_WIRE_1 : _ar_ready_WIRE_0; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_2 = Queue_2_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_2 = 6'h2 == auto_in_ar_bits_id ? _ar_ready_WIRE_2 : _GEN_1; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_3 = Queue_3_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_3 = 6'h3 == auto_in_ar_bits_id ? _ar_ready_WIRE_3 : _GEN_2; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_4 = Queue_4_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_4 = 6'h4 == auto_in_ar_bits_id ? _ar_ready_WIRE_4 : _GEN_3; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_5 = Queue_5_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_5 = 6'h5 == auto_in_ar_bits_id ? _ar_ready_WIRE_5 : _GEN_4; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_6 = Queue_6_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_6 = 6'h6 == auto_in_ar_bits_id ? _ar_ready_WIRE_6 : _GEN_5; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_7 = Queue_7_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_7 = 6'h7 == auto_in_ar_bits_id ? _ar_ready_WIRE_7 : _GEN_6; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_8 = Queue_8_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_8 = 6'h8 == auto_in_ar_bits_id ? _ar_ready_WIRE_8 : _GEN_7; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_9 = Queue_9_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_9 = 6'h9 == auto_in_ar_bits_id ? _ar_ready_WIRE_9 : _GEN_8; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_10 = Queue_10_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_10 = 6'ha == auto_in_ar_bits_id ? _ar_ready_WIRE_10 : _GEN_9; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_11 = Queue_11_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_11 = 6'hb == auto_in_ar_bits_id ? _ar_ready_WIRE_11 : _GEN_10; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_12 = Queue_12_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_12 = 6'hc == auto_in_ar_bits_id ? _ar_ready_WIRE_12 : _GEN_11; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_13 = Queue_13_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_13 = 6'hd == auto_in_ar_bits_id ? _ar_ready_WIRE_13 : _GEN_12; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_14 = Queue_14_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_14 = 6'he == auto_in_ar_bits_id ? _ar_ready_WIRE_14 : _GEN_13; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_15 = Queue_15_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_15 = 6'hf == auto_in_ar_bits_id ? _ar_ready_WIRE_15 : _GEN_14; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_16 = Queue_16_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_16 = 6'h10 == auto_in_ar_bits_id ? _ar_ready_WIRE_16 : _GEN_15; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_17 = Queue_17_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_17 = 6'h11 == auto_in_ar_bits_id ? _ar_ready_WIRE_17 : _GEN_16; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_18 = Queue_18_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_18 = 6'h12 == auto_in_ar_bits_id ? _ar_ready_WIRE_18 : _GEN_17; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_19 = Queue_19_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_19 = 6'h13 == auto_in_ar_bits_id ? _ar_ready_WIRE_19 : _GEN_18; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_20 = Queue_20_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_20 = 6'h14 == auto_in_ar_bits_id ? _ar_ready_WIRE_20 : _GEN_19; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_21 = Queue_21_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_21 = 6'h15 == auto_in_ar_bits_id ? _ar_ready_WIRE_21 : _GEN_20; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_22 = Queue_22_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_22 = 6'h16 == auto_in_ar_bits_id ? _ar_ready_WIRE_22 : _GEN_21; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_23 = Queue_23_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_23 = 6'h17 == auto_in_ar_bits_id ? _ar_ready_WIRE_23 : _GEN_22; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_24 = Queue_24_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_24 = 6'h18 == auto_in_ar_bits_id ? _ar_ready_WIRE_24 : _GEN_23; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_25 = Queue_25_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_25 = 6'h19 == auto_in_ar_bits_id ? _ar_ready_WIRE_25 : _GEN_24; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_26 = Queue_26_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_26 = 6'h1a == auto_in_ar_bits_id ? _ar_ready_WIRE_26 : _GEN_25; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_27 = Queue_27_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_27 = 6'h1b == auto_in_ar_bits_id ? _ar_ready_WIRE_27 : _GEN_26; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_28 = Queue_28_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_28 = 6'h1c == auto_in_ar_bits_id ? _ar_ready_WIRE_28 : _GEN_27; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_29 = Queue_29_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_29 = 6'h1d == auto_in_ar_bits_id ? _ar_ready_WIRE_29 : _GEN_28; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_30 = Queue_30_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_30 = 6'h1e == auto_in_ar_bits_id ? _ar_ready_WIRE_30 : _GEN_29; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_31 = Queue_31_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_31 = 6'h1f == auto_in_ar_bits_id ? _ar_ready_WIRE_31 : _GEN_30; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_32 = Queue_32_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_32 = 6'h20 == auto_in_ar_bits_id ? _ar_ready_WIRE_32 : _GEN_31; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_33 = Queue_33_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_33 = 6'h21 == auto_in_ar_bits_id ? _ar_ready_WIRE_33 : _GEN_32; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_34 = Queue_34_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_34 = 6'h22 == auto_in_ar_bits_id ? _ar_ready_WIRE_34 : _GEN_33; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_35 = Queue_35_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_35 = 6'h23 == auto_in_ar_bits_id ? _ar_ready_WIRE_35 : _GEN_34; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_36 = Queue_36_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_36 = 6'h24 == auto_in_ar_bits_id ? _ar_ready_WIRE_36 : _GEN_35; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_37 = Queue_37_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_37 = 6'h25 == auto_in_ar_bits_id ? _ar_ready_WIRE_37 : _GEN_36; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_38 = Queue_38_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_38 = 6'h26 == auto_in_ar_bits_id ? _ar_ready_WIRE_38 : _GEN_37; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_39 = Queue_39_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_39 = 6'h27 == auto_in_ar_bits_id ? _ar_ready_WIRE_39 : _GEN_38; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_40 = Queue_40_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_40 = 6'h28 == auto_in_ar_bits_id ? _ar_ready_WIRE_40 : _GEN_39; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_41 = Queue_41_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_41 = 6'h29 == auto_in_ar_bits_id ? _ar_ready_WIRE_41 : _GEN_40; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_42 = Queue_42_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_42 = 6'h2a == auto_in_ar_bits_id ? _ar_ready_WIRE_42 : _GEN_41; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_43 = Queue_43_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_43 = 6'h2b == auto_in_ar_bits_id ? _ar_ready_WIRE_43 : _GEN_42; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_44 = Queue_44_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_44 = 6'h2c == auto_in_ar_bits_id ? _ar_ready_WIRE_44 : _GEN_43; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_45 = Queue_45_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_45 = 6'h2d == auto_in_ar_bits_id ? _ar_ready_WIRE_45 : _GEN_44; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_46 = Queue_46_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_46 = 6'h2e == auto_in_ar_bits_id ? _ar_ready_WIRE_46 : _GEN_45; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_47 = Queue_47_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_47 = 6'h2f == auto_in_ar_bits_id ? _ar_ready_WIRE_47 : _GEN_46; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_48 = Queue_48_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_48 = 6'h30 == auto_in_ar_bits_id ? _ar_ready_WIRE_48 : _GEN_47; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_49 = Queue_49_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_49 = 6'h31 == auto_in_ar_bits_id ? _ar_ready_WIRE_49 : _GEN_48; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_50 = Queue_50_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_50 = 6'h32 == auto_in_ar_bits_id ? _ar_ready_WIRE_50 : _GEN_49; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_51 = Queue_51_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_51 = 6'h33 == auto_in_ar_bits_id ? _ar_ready_WIRE_51 : _GEN_50; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_52 = Queue_52_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_52 = 6'h34 == auto_in_ar_bits_id ? _ar_ready_WIRE_52 : _GEN_51; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_53 = Queue_53_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_53 = 6'h35 == auto_in_ar_bits_id ? _ar_ready_WIRE_53 : _GEN_52; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_54 = Queue_54_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_54 = 6'h36 == auto_in_ar_bits_id ? _ar_ready_WIRE_54 : _GEN_53; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_55 = Queue_55_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_55 = 6'h37 == auto_in_ar_bits_id ? _ar_ready_WIRE_55 : _GEN_54; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_56 = Queue_56_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_56 = 6'h38 == auto_in_ar_bits_id ? _ar_ready_WIRE_56 : _GEN_55; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_57 = Queue_57_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_57 = 6'h39 == auto_in_ar_bits_id ? _ar_ready_WIRE_57 : _GEN_56; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_58 = Queue_58_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_58 = 6'h3a == auto_in_ar_bits_id ? _ar_ready_WIRE_58 : _GEN_57; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_59 = Queue_59_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_59 = 6'h3b == auto_in_ar_bits_id ? _ar_ready_WIRE_59 : _GEN_58; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_60 = Queue_60_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_60 = 6'h3c == auto_in_ar_bits_id ? _ar_ready_WIRE_60 : _GEN_59; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_61 = Queue_61_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_61 = 6'h3d == auto_in_ar_bits_id ? _ar_ready_WIRE_61 : _GEN_60; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_62 = Queue_62_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_62 = 6'h3e == auto_in_ar_bits_id ? _ar_ready_WIRE_62 : _GEN_61; // @[UserYanker.scala 59:{36,36}]
  wire  _ar_ready_WIRE_63 = Queue_63_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_63 = 6'h3f == auto_in_ar_bits_id ? _ar_ready_WIRE_63 : _GEN_62; // @[UserYanker.scala 59:{36,36}]
  wire  _r_valid_WIRE_0 = Queue_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _r_valid_WIRE_1 = Queue_1_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_65 = 6'h1 == auto_out_r_bits_id ? _r_valid_WIRE_1 : _r_valid_WIRE_0; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_2 = Queue_2_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_66 = 6'h2 == auto_out_r_bits_id ? _r_valid_WIRE_2 : _GEN_65; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_3 = Queue_3_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_67 = 6'h3 == auto_out_r_bits_id ? _r_valid_WIRE_3 : _GEN_66; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_4 = Queue_4_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_68 = 6'h4 == auto_out_r_bits_id ? _r_valid_WIRE_4 : _GEN_67; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_5 = Queue_5_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_69 = 6'h5 == auto_out_r_bits_id ? _r_valid_WIRE_5 : _GEN_68; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_6 = Queue_6_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_70 = 6'h6 == auto_out_r_bits_id ? _r_valid_WIRE_6 : _GEN_69; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_7 = Queue_7_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_71 = 6'h7 == auto_out_r_bits_id ? _r_valid_WIRE_7 : _GEN_70; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_8 = Queue_8_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_72 = 6'h8 == auto_out_r_bits_id ? _r_valid_WIRE_8 : _GEN_71; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_9 = Queue_9_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_73 = 6'h9 == auto_out_r_bits_id ? _r_valid_WIRE_9 : _GEN_72; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_10 = Queue_10_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_74 = 6'ha == auto_out_r_bits_id ? _r_valid_WIRE_10 : _GEN_73; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_11 = Queue_11_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_75 = 6'hb == auto_out_r_bits_id ? _r_valid_WIRE_11 : _GEN_74; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_12 = Queue_12_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_76 = 6'hc == auto_out_r_bits_id ? _r_valid_WIRE_12 : _GEN_75; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_13 = Queue_13_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_77 = 6'hd == auto_out_r_bits_id ? _r_valid_WIRE_13 : _GEN_76; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_14 = Queue_14_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_78 = 6'he == auto_out_r_bits_id ? _r_valid_WIRE_14 : _GEN_77; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_15 = Queue_15_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_79 = 6'hf == auto_out_r_bits_id ? _r_valid_WIRE_15 : _GEN_78; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_16 = Queue_16_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_80 = 6'h10 == auto_out_r_bits_id ? _r_valid_WIRE_16 : _GEN_79; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_17 = Queue_17_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_81 = 6'h11 == auto_out_r_bits_id ? _r_valid_WIRE_17 : _GEN_80; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_18 = Queue_18_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_82 = 6'h12 == auto_out_r_bits_id ? _r_valid_WIRE_18 : _GEN_81; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_19 = Queue_19_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_83 = 6'h13 == auto_out_r_bits_id ? _r_valid_WIRE_19 : _GEN_82; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_20 = Queue_20_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_84 = 6'h14 == auto_out_r_bits_id ? _r_valid_WIRE_20 : _GEN_83; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_21 = Queue_21_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_85 = 6'h15 == auto_out_r_bits_id ? _r_valid_WIRE_21 : _GEN_84; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_22 = Queue_22_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_86 = 6'h16 == auto_out_r_bits_id ? _r_valid_WIRE_22 : _GEN_85; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_23 = Queue_23_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_87 = 6'h17 == auto_out_r_bits_id ? _r_valid_WIRE_23 : _GEN_86; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_24 = Queue_24_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_88 = 6'h18 == auto_out_r_bits_id ? _r_valid_WIRE_24 : _GEN_87; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_25 = Queue_25_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_89 = 6'h19 == auto_out_r_bits_id ? _r_valid_WIRE_25 : _GEN_88; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_26 = Queue_26_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_90 = 6'h1a == auto_out_r_bits_id ? _r_valid_WIRE_26 : _GEN_89; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_27 = Queue_27_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_91 = 6'h1b == auto_out_r_bits_id ? _r_valid_WIRE_27 : _GEN_90; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_28 = Queue_28_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_92 = 6'h1c == auto_out_r_bits_id ? _r_valid_WIRE_28 : _GEN_91; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_29 = Queue_29_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_93 = 6'h1d == auto_out_r_bits_id ? _r_valid_WIRE_29 : _GEN_92; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_30 = Queue_30_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_94 = 6'h1e == auto_out_r_bits_id ? _r_valid_WIRE_30 : _GEN_93; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_31 = Queue_31_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_95 = 6'h1f == auto_out_r_bits_id ? _r_valid_WIRE_31 : _GEN_94; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_32 = Queue_32_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_96 = 6'h20 == auto_out_r_bits_id ? _r_valid_WIRE_32 : _GEN_95; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_33 = Queue_33_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_97 = 6'h21 == auto_out_r_bits_id ? _r_valid_WIRE_33 : _GEN_96; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_34 = Queue_34_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_98 = 6'h22 == auto_out_r_bits_id ? _r_valid_WIRE_34 : _GEN_97; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_35 = Queue_35_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_99 = 6'h23 == auto_out_r_bits_id ? _r_valid_WIRE_35 : _GEN_98; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_36 = Queue_36_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_100 = 6'h24 == auto_out_r_bits_id ? _r_valid_WIRE_36 : _GEN_99; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_37 = Queue_37_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_101 = 6'h25 == auto_out_r_bits_id ? _r_valid_WIRE_37 : _GEN_100; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_38 = Queue_38_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_102 = 6'h26 == auto_out_r_bits_id ? _r_valid_WIRE_38 : _GEN_101; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_39 = Queue_39_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_103 = 6'h27 == auto_out_r_bits_id ? _r_valid_WIRE_39 : _GEN_102; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_40 = Queue_40_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_104 = 6'h28 == auto_out_r_bits_id ? _r_valid_WIRE_40 : _GEN_103; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_41 = Queue_41_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_105 = 6'h29 == auto_out_r_bits_id ? _r_valid_WIRE_41 : _GEN_104; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_42 = Queue_42_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_106 = 6'h2a == auto_out_r_bits_id ? _r_valid_WIRE_42 : _GEN_105; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_43 = Queue_43_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_107 = 6'h2b == auto_out_r_bits_id ? _r_valid_WIRE_43 : _GEN_106; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_44 = Queue_44_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_108 = 6'h2c == auto_out_r_bits_id ? _r_valid_WIRE_44 : _GEN_107; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_45 = Queue_45_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_109 = 6'h2d == auto_out_r_bits_id ? _r_valid_WIRE_45 : _GEN_108; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_46 = Queue_46_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_110 = 6'h2e == auto_out_r_bits_id ? _r_valid_WIRE_46 : _GEN_109; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_47 = Queue_47_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_111 = 6'h2f == auto_out_r_bits_id ? _r_valid_WIRE_47 : _GEN_110; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_48 = Queue_48_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_112 = 6'h30 == auto_out_r_bits_id ? _r_valid_WIRE_48 : _GEN_111; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_49 = Queue_49_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_113 = 6'h31 == auto_out_r_bits_id ? _r_valid_WIRE_49 : _GEN_112; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_50 = Queue_50_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_114 = 6'h32 == auto_out_r_bits_id ? _r_valid_WIRE_50 : _GEN_113; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_51 = Queue_51_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_115 = 6'h33 == auto_out_r_bits_id ? _r_valid_WIRE_51 : _GEN_114; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_52 = Queue_52_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_116 = 6'h34 == auto_out_r_bits_id ? _r_valid_WIRE_52 : _GEN_115; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_53 = Queue_53_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_117 = 6'h35 == auto_out_r_bits_id ? _r_valid_WIRE_53 : _GEN_116; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_54 = Queue_54_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_118 = 6'h36 == auto_out_r_bits_id ? _r_valid_WIRE_54 : _GEN_117; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_55 = Queue_55_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_119 = 6'h37 == auto_out_r_bits_id ? _r_valid_WIRE_55 : _GEN_118; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_56 = Queue_56_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_120 = 6'h38 == auto_out_r_bits_id ? _r_valid_WIRE_56 : _GEN_119; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_57 = Queue_57_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_121 = 6'h39 == auto_out_r_bits_id ? _r_valid_WIRE_57 : _GEN_120; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_58 = Queue_58_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_122 = 6'h3a == auto_out_r_bits_id ? _r_valid_WIRE_58 : _GEN_121; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_59 = Queue_59_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_123 = 6'h3b == auto_out_r_bits_id ? _r_valid_WIRE_59 : _GEN_122; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_60 = Queue_60_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_124 = 6'h3c == auto_out_r_bits_id ? _r_valid_WIRE_60 : _GEN_123; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_61 = Queue_61_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_125 = 6'h3d == auto_out_r_bits_id ? _r_valid_WIRE_61 : _GEN_124; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_62 = Queue_62_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_126 = 6'h3e == auto_out_r_bits_id ? _r_valid_WIRE_62 : _GEN_125; // @[UserYanker.scala 66:{28,28}]
  wire  _r_valid_WIRE_63 = Queue_63_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_127 = 6'h3f == auto_out_r_bits_id ? _r_valid_WIRE_63 : _GEN_126; // @[UserYanker.scala 66:{28,28}]
  wire  _T_3 = ~reset; // @[UserYanker.scala 66:14]
  wire [1:0] _r_bits_WIRE_0_extra_id = Queue_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _r_bits_WIRE_1_extra_id = Queue_1_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_129 = 6'h1 == auto_out_r_bits_id ? _r_bits_WIRE_1_extra_id : _r_bits_WIRE_0_extra_id; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_2_extra_id = Queue_2_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_130 = 6'h2 == auto_out_r_bits_id ? _r_bits_WIRE_2_extra_id : _GEN_129; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_3_extra_id = Queue_3_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_131 = 6'h3 == auto_out_r_bits_id ? _r_bits_WIRE_3_extra_id : _GEN_130; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_4_extra_id = Queue_4_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_132 = 6'h4 == auto_out_r_bits_id ? _r_bits_WIRE_4_extra_id : _GEN_131; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_5_extra_id = Queue_5_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_133 = 6'h5 == auto_out_r_bits_id ? _r_bits_WIRE_5_extra_id : _GEN_132; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_6_extra_id = Queue_6_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_134 = 6'h6 == auto_out_r_bits_id ? _r_bits_WIRE_6_extra_id : _GEN_133; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_7_extra_id = Queue_7_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_135 = 6'h7 == auto_out_r_bits_id ? _r_bits_WIRE_7_extra_id : _GEN_134; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_8_extra_id = Queue_8_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_136 = 6'h8 == auto_out_r_bits_id ? _r_bits_WIRE_8_extra_id : _GEN_135; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_9_extra_id = Queue_9_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_137 = 6'h9 == auto_out_r_bits_id ? _r_bits_WIRE_9_extra_id : _GEN_136; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_10_extra_id = Queue_10_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_138 = 6'ha == auto_out_r_bits_id ? _r_bits_WIRE_10_extra_id : _GEN_137; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_11_extra_id = Queue_11_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_139 = 6'hb == auto_out_r_bits_id ? _r_bits_WIRE_11_extra_id : _GEN_138; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_12_extra_id = Queue_12_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_140 = 6'hc == auto_out_r_bits_id ? _r_bits_WIRE_12_extra_id : _GEN_139; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_13_extra_id = Queue_13_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_141 = 6'hd == auto_out_r_bits_id ? _r_bits_WIRE_13_extra_id : _GEN_140; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_14_extra_id = Queue_14_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_142 = 6'he == auto_out_r_bits_id ? _r_bits_WIRE_14_extra_id : _GEN_141; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_15_extra_id = Queue_15_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_143 = 6'hf == auto_out_r_bits_id ? _r_bits_WIRE_15_extra_id : _GEN_142; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_16_extra_id = Queue_16_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_144 = 6'h10 == auto_out_r_bits_id ? _r_bits_WIRE_16_extra_id : _GEN_143; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_17_extra_id = Queue_17_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_145 = 6'h11 == auto_out_r_bits_id ? _r_bits_WIRE_17_extra_id : _GEN_144; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_18_extra_id = Queue_18_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_146 = 6'h12 == auto_out_r_bits_id ? _r_bits_WIRE_18_extra_id : _GEN_145; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_19_extra_id = Queue_19_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_147 = 6'h13 == auto_out_r_bits_id ? _r_bits_WIRE_19_extra_id : _GEN_146; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_20_extra_id = Queue_20_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_148 = 6'h14 == auto_out_r_bits_id ? _r_bits_WIRE_20_extra_id : _GEN_147; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_21_extra_id = Queue_21_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_149 = 6'h15 == auto_out_r_bits_id ? _r_bits_WIRE_21_extra_id : _GEN_148; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_22_extra_id = Queue_22_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_150 = 6'h16 == auto_out_r_bits_id ? _r_bits_WIRE_22_extra_id : _GEN_149; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_23_extra_id = Queue_23_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_151 = 6'h17 == auto_out_r_bits_id ? _r_bits_WIRE_23_extra_id : _GEN_150; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_24_extra_id = Queue_24_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_152 = 6'h18 == auto_out_r_bits_id ? _r_bits_WIRE_24_extra_id : _GEN_151; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_25_extra_id = Queue_25_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_153 = 6'h19 == auto_out_r_bits_id ? _r_bits_WIRE_25_extra_id : _GEN_152; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_26_extra_id = Queue_26_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_154 = 6'h1a == auto_out_r_bits_id ? _r_bits_WIRE_26_extra_id : _GEN_153; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_27_extra_id = Queue_27_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_155 = 6'h1b == auto_out_r_bits_id ? _r_bits_WIRE_27_extra_id : _GEN_154; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_28_extra_id = Queue_28_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_156 = 6'h1c == auto_out_r_bits_id ? _r_bits_WIRE_28_extra_id : _GEN_155; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_29_extra_id = Queue_29_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_157 = 6'h1d == auto_out_r_bits_id ? _r_bits_WIRE_29_extra_id : _GEN_156; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_30_extra_id = Queue_30_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_158 = 6'h1e == auto_out_r_bits_id ? _r_bits_WIRE_30_extra_id : _GEN_157; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_31_extra_id = Queue_31_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_159 = 6'h1f == auto_out_r_bits_id ? _r_bits_WIRE_31_extra_id : _GEN_158; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_32_extra_id = Queue_32_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_160 = 6'h20 == auto_out_r_bits_id ? _r_bits_WIRE_32_extra_id : _GEN_159; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_33_extra_id = Queue_33_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_161 = 6'h21 == auto_out_r_bits_id ? _r_bits_WIRE_33_extra_id : _GEN_160; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_34_extra_id = Queue_34_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_162 = 6'h22 == auto_out_r_bits_id ? _r_bits_WIRE_34_extra_id : _GEN_161; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_35_extra_id = Queue_35_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_163 = 6'h23 == auto_out_r_bits_id ? _r_bits_WIRE_35_extra_id : _GEN_162; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_36_extra_id = Queue_36_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_164 = 6'h24 == auto_out_r_bits_id ? _r_bits_WIRE_36_extra_id : _GEN_163; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_37_extra_id = Queue_37_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_165 = 6'h25 == auto_out_r_bits_id ? _r_bits_WIRE_37_extra_id : _GEN_164; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_38_extra_id = Queue_38_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_166 = 6'h26 == auto_out_r_bits_id ? _r_bits_WIRE_38_extra_id : _GEN_165; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_39_extra_id = Queue_39_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_167 = 6'h27 == auto_out_r_bits_id ? _r_bits_WIRE_39_extra_id : _GEN_166; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_40_extra_id = Queue_40_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_168 = 6'h28 == auto_out_r_bits_id ? _r_bits_WIRE_40_extra_id : _GEN_167; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_41_extra_id = Queue_41_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_169 = 6'h29 == auto_out_r_bits_id ? _r_bits_WIRE_41_extra_id : _GEN_168; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_42_extra_id = Queue_42_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_170 = 6'h2a == auto_out_r_bits_id ? _r_bits_WIRE_42_extra_id : _GEN_169; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_43_extra_id = Queue_43_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_171 = 6'h2b == auto_out_r_bits_id ? _r_bits_WIRE_43_extra_id : _GEN_170; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_44_extra_id = Queue_44_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_172 = 6'h2c == auto_out_r_bits_id ? _r_bits_WIRE_44_extra_id : _GEN_171; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_45_extra_id = Queue_45_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_173 = 6'h2d == auto_out_r_bits_id ? _r_bits_WIRE_45_extra_id : _GEN_172; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_46_extra_id = Queue_46_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_174 = 6'h2e == auto_out_r_bits_id ? _r_bits_WIRE_46_extra_id : _GEN_173; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_47_extra_id = Queue_47_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_175 = 6'h2f == auto_out_r_bits_id ? _r_bits_WIRE_47_extra_id : _GEN_174; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_48_extra_id = Queue_48_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_176 = 6'h30 == auto_out_r_bits_id ? _r_bits_WIRE_48_extra_id : _GEN_175; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_49_extra_id = Queue_49_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_177 = 6'h31 == auto_out_r_bits_id ? _r_bits_WIRE_49_extra_id : _GEN_176; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_50_extra_id = Queue_50_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_178 = 6'h32 == auto_out_r_bits_id ? _r_bits_WIRE_50_extra_id : _GEN_177; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_51_extra_id = Queue_51_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_179 = 6'h33 == auto_out_r_bits_id ? _r_bits_WIRE_51_extra_id : _GEN_178; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_52_extra_id = Queue_52_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_180 = 6'h34 == auto_out_r_bits_id ? _r_bits_WIRE_52_extra_id : _GEN_179; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_53_extra_id = Queue_53_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_181 = 6'h35 == auto_out_r_bits_id ? _r_bits_WIRE_53_extra_id : _GEN_180; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_54_extra_id = Queue_54_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_182 = 6'h36 == auto_out_r_bits_id ? _r_bits_WIRE_54_extra_id : _GEN_181; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_55_extra_id = Queue_55_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_183 = 6'h37 == auto_out_r_bits_id ? _r_bits_WIRE_55_extra_id : _GEN_182; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_56_extra_id = Queue_56_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_184 = 6'h38 == auto_out_r_bits_id ? _r_bits_WIRE_56_extra_id : _GEN_183; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_57_extra_id = Queue_57_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_185 = 6'h39 == auto_out_r_bits_id ? _r_bits_WIRE_57_extra_id : _GEN_184; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_58_extra_id = Queue_58_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_186 = 6'h3a == auto_out_r_bits_id ? _r_bits_WIRE_58_extra_id : _GEN_185; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_59_extra_id = Queue_59_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_187 = 6'h3b == auto_out_r_bits_id ? _r_bits_WIRE_59_extra_id : _GEN_186; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_60_extra_id = Queue_60_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_188 = 6'h3c == auto_out_r_bits_id ? _r_bits_WIRE_60_extra_id : _GEN_187; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_61_extra_id = Queue_61_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_189 = 6'h3d == auto_out_r_bits_id ? _r_bits_WIRE_61_extra_id : _GEN_188; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_62_extra_id = Queue_62_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _GEN_190 = 6'h3e == auto_out_r_bits_id ? _r_bits_WIRE_62_extra_id : _GEN_189; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _r_bits_WIRE_63_extra_id = Queue_63_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _r_bits_WIRE_0_tl_state_source = Queue_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _r_bits_WIRE_1_tl_state_source = Queue_1_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_193 = 6'h1 == auto_out_r_bits_id ? _r_bits_WIRE_1_tl_state_source : _r_bits_WIRE_0_tl_state_source; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_2_tl_state_source = Queue_2_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_194 = 6'h2 == auto_out_r_bits_id ? _r_bits_WIRE_2_tl_state_source : _GEN_193; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_3_tl_state_source = Queue_3_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_195 = 6'h3 == auto_out_r_bits_id ? _r_bits_WIRE_3_tl_state_source : _GEN_194; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_4_tl_state_source = Queue_4_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_196 = 6'h4 == auto_out_r_bits_id ? _r_bits_WIRE_4_tl_state_source : _GEN_195; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_5_tl_state_source = Queue_5_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_197 = 6'h5 == auto_out_r_bits_id ? _r_bits_WIRE_5_tl_state_source : _GEN_196; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_6_tl_state_source = Queue_6_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_198 = 6'h6 == auto_out_r_bits_id ? _r_bits_WIRE_6_tl_state_source : _GEN_197; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_7_tl_state_source = Queue_7_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_199 = 6'h7 == auto_out_r_bits_id ? _r_bits_WIRE_7_tl_state_source : _GEN_198; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_8_tl_state_source = Queue_8_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_200 = 6'h8 == auto_out_r_bits_id ? _r_bits_WIRE_8_tl_state_source : _GEN_199; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_9_tl_state_source = Queue_9_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_201 = 6'h9 == auto_out_r_bits_id ? _r_bits_WIRE_9_tl_state_source : _GEN_200; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_10_tl_state_source = Queue_10_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_202 = 6'ha == auto_out_r_bits_id ? _r_bits_WIRE_10_tl_state_source : _GEN_201; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_11_tl_state_source = Queue_11_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_203 = 6'hb == auto_out_r_bits_id ? _r_bits_WIRE_11_tl_state_source : _GEN_202; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_12_tl_state_source = Queue_12_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_204 = 6'hc == auto_out_r_bits_id ? _r_bits_WIRE_12_tl_state_source : _GEN_203; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_13_tl_state_source = Queue_13_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_205 = 6'hd == auto_out_r_bits_id ? _r_bits_WIRE_13_tl_state_source : _GEN_204; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_14_tl_state_source = Queue_14_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_206 = 6'he == auto_out_r_bits_id ? _r_bits_WIRE_14_tl_state_source : _GEN_205; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_15_tl_state_source = Queue_15_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_207 = 6'hf == auto_out_r_bits_id ? _r_bits_WIRE_15_tl_state_source : _GEN_206; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_16_tl_state_source = Queue_16_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_208 = 6'h10 == auto_out_r_bits_id ? _r_bits_WIRE_16_tl_state_source : _GEN_207; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_17_tl_state_source = Queue_17_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_209 = 6'h11 == auto_out_r_bits_id ? _r_bits_WIRE_17_tl_state_source : _GEN_208; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_18_tl_state_source = Queue_18_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_210 = 6'h12 == auto_out_r_bits_id ? _r_bits_WIRE_18_tl_state_source : _GEN_209; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_19_tl_state_source = Queue_19_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_211 = 6'h13 == auto_out_r_bits_id ? _r_bits_WIRE_19_tl_state_source : _GEN_210; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_20_tl_state_source = Queue_20_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_212 = 6'h14 == auto_out_r_bits_id ? _r_bits_WIRE_20_tl_state_source : _GEN_211; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_21_tl_state_source = Queue_21_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_213 = 6'h15 == auto_out_r_bits_id ? _r_bits_WIRE_21_tl_state_source : _GEN_212; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_22_tl_state_source = Queue_22_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_214 = 6'h16 == auto_out_r_bits_id ? _r_bits_WIRE_22_tl_state_source : _GEN_213; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_23_tl_state_source = Queue_23_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_215 = 6'h17 == auto_out_r_bits_id ? _r_bits_WIRE_23_tl_state_source : _GEN_214; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_24_tl_state_source = Queue_24_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_216 = 6'h18 == auto_out_r_bits_id ? _r_bits_WIRE_24_tl_state_source : _GEN_215; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_25_tl_state_source = Queue_25_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_217 = 6'h19 == auto_out_r_bits_id ? _r_bits_WIRE_25_tl_state_source : _GEN_216; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_26_tl_state_source = Queue_26_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_218 = 6'h1a == auto_out_r_bits_id ? _r_bits_WIRE_26_tl_state_source : _GEN_217; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_27_tl_state_source = Queue_27_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_219 = 6'h1b == auto_out_r_bits_id ? _r_bits_WIRE_27_tl_state_source : _GEN_218; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_28_tl_state_source = Queue_28_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_220 = 6'h1c == auto_out_r_bits_id ? _r_bits_WIRE_28_tl_state_source : _GEN_219; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_29_tl_state_source = Queue_29_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_221 = 6'h1d == auto_out_r_bits_id ? _r_bits_WIRE_29_tl_state_source : _GEN_220; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_30_tl_state_source = Queue_30_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_222 = 6'h1e == auto_out_r_bits_id ? _r_bits_WIRE_30_tl_state_source : _GEN_221; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_31_tl_state_source = Queue_31_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_223 = 6'h1f == auto_out_r_bits_id ? _r_bits_WIRE_31_tl_state_source : _GEN_222; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_32_tl_state_source = Queue_32_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_224 = 6'h20 == auto_out_r_bits_id ? _r_bits_WIRE_32_tl_state_source : _GEN_223; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_33_tl_state_source = Queue_33_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_225 = 6'h21 == auto_out_r_bits_id ? _r_bits_WIRE_33_tl_state_source : _GEN_224; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_34_tl_state_source = Queue_34_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_226 = 6'h22 == auto_out_r_bits_id ? _r_bits_WIRE_34_tl_state_source : _GEN_225; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_35_tl_state_source = Queue_35_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_227 = 6'h23 == auto_out_r_bits_id ? _r_bits_WIRE_35_tl_state_source : _GEN_226; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_36_tl_state_source = Queue_36_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_228 = 6'h24 == auto_out_r_bits_id ? _r_bits_WIRE_36_tl_state_source : _GEN_227; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_37_tl_state_source = Queue_37_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_229 = 6'h25 == auto_out_r_bits_id ? _r_bits_WIRE_37_tl_state_source : _GEN_228; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_38_tl_state_source = Queue_38_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_230 = 6'h26 == auto_out_r_bits_id ? _r_bits_WIRE_38_tl_state_source : _GEN_229; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_39_tl_state_source = Queue_39_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_231 = 6'h27 == auto_out_r_bits_id ? _r_bits_WIRE_39_tl_state_source : _GEN_230; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_40_tl_state_source = Queue_40_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_232 = 6'h28 == auto_out_r_bits_id ? _r_bits_WIRE_40_tl_state_source : _GEN_231; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_41_tl_state_source = Queue_41_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_233 = 6'h29 == auto_out_r_bits_id ? _r_bits_WIRE_41_tl_state_source : _GEN_232; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_42_tl_state_source = Queue_42_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_234 = 6'h2a == auto_out_r_bits_id ? _r_bits_WIRE_42_tl_state_source : _GEN_233; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_43_tl_state_source = Queue_43_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_235 = 6'h2b == auto_out_r_bits_id ? _r_bits_WIRE_43_tl_state_source : _GEN_234; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_44_tl_state_source = Queue_44_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_236 = 6'h2c == auto_out_r_bits_id ? _r_bits_WIRE_44_tl_state_source : _GEN_235; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_45_tl_state_source = Queue_45_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_237 = 6'h2d == auto_out_r_bits_id ? _r_bits_WIRE_45_tl_state_source : _GEN_236; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_46_tl_state_source = Queue_46_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_238 = 6'h2e == auto_out_r_bits_id ? _r_bits_WIRE_46_tl_state_source : _GEN_237; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_47_tl_state_source = Queue_47_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_239 = 6'h2f == auto_out_r_bits_id ? _r_bits_WIRE_47_tl_state_source : _GEN_238; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_48_tl_state_source = Queue_48_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_240 = 6'h30 == auto_out_r_bits_id ? _r_bits_WIRE_48_tl_state_source : _GEN_239; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_49_tl_state_source = Queue_49_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_241 = 6'h31 == auto_out_r_bits_id ? _r_bits_WIRE_49_tl_state_source : _GEN_240; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_50_tl_state_source = Queue_50_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_242 = 6'h32 == auto_out_r_bits_id ? _r_bits_WIRE_50_tl_state_source : _GEN_241; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_51_tl_state_source = Queue_51_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_243 = 6'h33 == auto_out_r_bits_id ? _r_bits_WIRE_51_tl_state_source : _GEN_242; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_52_tl_state_source = Queue_52_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_244 = 6'h34 == auto_out_r_bits_id ? _r_bits_WIRE_52_tl_state_source : _GEN_243; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_53_tl_state_source = Queue_53_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_245 = 6'h35 == auto_out_r_bits_id ? _r_bits_WIRE_53_tl_state_source : _GEN_244; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_54_tl_state_source = Queue_54_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_246 = 6'h36 == auto_out_r_bits_id ? _r_bits_WIRE_54_tl_state_source : _GEN_245; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_55_tl_state_source = Queue_55_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_247 = 6'h37 == auto_out_r_bits_id ? _r_bits_WIRE_55_tl_state_source : _GEN_246; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_56_tl_state_source = Queue_56_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_248 = 6'h38 == auto_out_r_bits_id ? _r_bits_WIRE_56_tl_state_source : _GEN_247; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_57_tl_state_source = Queue_57_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_249 = 6'h39 == auto_out_r_bits_id ? _r_bits_WIRE_57_tl_state_source : _GEN_248; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_58_tl_state_source = Queue_58_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_250 = 6'h3a == auto_out_r_bits_id ? _r_bits_WIRE_58_tl_state_source : _GEN_249; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_59_tl_state_source = Queue_59_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_251 = 6'h3b == auto_out_r_bits_id ? _r_bits_WIRE_59_tl_state_source : _GEN_250; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_60_tl_state_source = Queue_60_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_252 = 6'h3c == auto_out_r_bits_id ? _r_bits_WIRE_60_tl_state_source : _GEN_251; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_61_tl_state_source = Queue_61_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_253 = 6'h3d == auto_out_r_bits_id ? _r_bits_WIRE_61_tl_state_source : _GEN_252; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_62_tl_state_source = Queue_62_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [6:0] _GEN_254 = 6'h3e == auto_out_r_bits_id ? _r_bits_WIRE_62_tl_state_source : _GEN_253; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _r_bits_WIRE_63_tl_state_source = Queue_63_io_deq_bits_tl_state_source; // @[UserYanker.scala 65:{27,27}]
  wire [63:0] _arsel_T = 64'h1 << auto_in_ar_bits_id; // @[OneHot.scala 64:12]
  wire  arsel_0 = _arsel_T[0]; // @[UserYanker.scala 70:55]
  wire  arsel_1 = _arsel_T[1]; // @[UserYanker.scala 70:55]
  wire  arsel_2 = _arsel_T[2]; // @[UserYanker.scala 70:55]
  wire  arsel_3 = _arsel_T[3]; // @[UserYanker.scala 70:55]
  wire  arsel_4 = _arsel_T[4]; // @[UserYanker.scala 70:55]
  wire  arsel_5 = _arsel_T[5]; // @[UserYanker.scala 70:55]
  wire  arsel_6 = _arsel_T[6]; // @[UserYanker.scala 70:55]
  wire  arsel_7 = _arsel_T[7]; // @[UserYanker.scala 70:55]
  wire  arsel_8 = _arsel_T[8]; // @[UserYanker.scala 70:55]
  wire  arsel_9 = _arsel_T[9]; // @[UserYanker.scala 70:55]
  wire  arsel_10 = _arsel_T[10]; // @[UserYanker.scala 70:55]
  wire  arsel_11 = _arsel_T[11]; // @[UserYanker.scala 70:55]
  wire  arsel_12 = _arsel_T[12]; // @[UserYanker.scala 70:55]
  wire  arsel_13 = _arsel_T[13]; // @[UserYanker.scala 70:55]
  wire  arsel_14 = _arsel_T[14]; // @[UserYanker.scala 70:55]
  wire  arsel_15 = _arsel_T[15]; // @[UserYanker.scala 70:55]
  wire  arsel_16 = _arsel_T[16]; // @[UserYanker.scala 70:55]
  wire  arsel_17 = _arsel_T[17]; // @[UserYanker.scala 70:55]
  wire  arsel_18 = _arsel_T[18]; // @[UserYanker.scala 70:55]
  wire  arsel_19 = _arsel_T[19]; // @[UserYanker.scala 70:55]
  wire  arsel_20 = _arsel_T[20]; // @[UserYanker.scala 70:55]
  wire  arsel_21 = _arsel_T[21]; // @[UserYanker.scala 70:55]
  wire  arsel_22 = _arsel_T[22]; // @[UserYanker.scala 70:55]
  wire  arsel_23 = _arsel_T[23]; // @[UserYanker.scala 70:55]
  wire  arsel_24 = _arsel_T[24]; // @[UserYanker.scala 70:55]
  wire  arsel_25 = _arsel_T[25]; // @[UserYanker.scala 70:55]
  wire  arsel_26 = _arsel_T[26]; // @[UserYanker.scala 70:55]
  wire  arsel_27 = _arsel_T[27]; // @[UserYanker.scala 70:55]
  wire  arsel_28 = _arsel_T[28]; // @[UserYanker.scala 70:55]
  wire  arsel_29 = _arsel_T[29]; // @[UserYanker.scala 70:55]
  wire  arsel_30 = _arsel_T[30]; // @[UserYanker.scala 70:55]
  wire  arsel_31 = _arsel_T[31]; // @[UserYanker.scala 70:55]
  wire  arsel_32 = _arsel_T[32]; // @[UserYanker.scala 70:55]
  wire  arsel_33 = _arsel_T[33]; // @[UserYanker.scala 70:55]
  wire  arsel_34 = _arsel_T[34]; // @[UserYanker.scala 70:55]
  wire  arsel_35 = _arsel_T[35]; // @[UserYanker.scala 70:55]
  wire  arsel_36 = _arsel_T[36]; // @[UserYanker.scala 70:55]
  wire  arsel_37 = _arsel_T[37]; // @[UserYanker.scala 70:55]
  wire  arsel_38 = _arsel_T[38]; // @[UserYanker.scala 70:55]
  wire  arsel_39 = _arsel_T[39]; // @[UserYanker.scala 70:55]
  wire  arsel_40 = _arsel_T[40]; // @[UserYanker.scala 70:55]
  wire  arsel_41 = _arsel_T[41]; // @[UserYanker.scala 70:55]
  wire  arsel_42 = _arsel_T[42]; // @[UserYanker.scala 70:55]
  wire  arsel_43 = _arsel_T[43]; // @[UserYanker.scala 70:55]
  wire  arsel_44 = _arsel_T[44]; // @[UserYanker.scala 70:55]
  wire  arsel_45 = _arsel_T[45]; // @[UserYanker.scala 70:55]
  wire  arsel_46 = _arsel_T[46]; // @[UserYanker.scala 70:55]
  wire  arsel_47 = _arsel_T[47]; // @[UserYanker.scala 70:55]
  wire  arsel_48 = _arsel_T[48]; // @[UserYanker.scala 70:55]
  wire  arsel_49 = _arsel_T[49]; // @[UserYanker.scala 70:55]
  wire  arsel_50 = _arsel_T[50]; // @[UserYanker.scala 70:55]
  wire  arsel_51 = _arsel_T[51]; // @[UserYanker.scala 70:55]
  wire  arsel_52 = _arsel_T[52]; // @[UserYanker.scala 70:55]
  wire  arsel_53 = _arsel_T[53]; // @[UserYanker.scala 70:55]
  wire  arsel_54 = _arsel_T[54]; // @[UserYanker.scala 70:55]
  wire  arsel_55 = _arsel_T[55]; // @[UserYanker.scala 70:55]
  wire  arsel_56 = _arsel_T[56]; // @[UserYanker.scala 70:55]
  wire  arsel_57 = _arsel_T[57]; // @[UserYanker.scala 70:55]
  wire  arsel_58 = _arsel_T[58]; // @[UserYanker.scala 70:55]
  wire  arsel_59 = _arsel_T[59]; // @[UserYanker.scala 70:55]
  wire  arsel_60 = _arsel_T[60]; // @[UserYanker.scala 70:55]
  wire  arsel_61 = _arsel_T[61]; // @[UserYanker.scala 70:55]
  wire  arsel_62 = _arsel_T[62]; // @[UserYanker.scala 70:55]
  wire  arsel_63 = _arsel_T[63]; // @[UserYanker.scala 70:55]
  wire [63:0] _rsel_T = 64'h1 << auto_out_r_bits_id; // @[OneHot.scala 64:12]
  wire  rsel_0 = _rsel_T[0]; // @[UserYanker.scala 71:55]
  wire  rsel_1 = _rsel_T[1]; // @[UserYanker.scala 71:55]
  wire  rsel_2 = _rsel_T[2]; // @[UserYanker.scala 71:55]
  wire  rsel_3 = _rsel_T[3]; // @[UserYanker.scala 71:55]
  wire  rsel_4 = _rsel_T[4]; // @[UserYanker.scala 71:55]
  wire  rsel_5 = _rsel_T[5]; // @[UserYanker.scala 71:55]
  wire  rsel_6 = _rsel_T[6]; // @[UserYanker.scala 71:55]
  wire  rsel_7 = _rsel_T[7]; // @[UserYanker.scala 71:55]
  wire  rsel_8 = _rsel_T[8]; // @[UserYanker.scala 71:55]
  wire  rsel_9 = _rsel_T[9]; // @[UserYanker.scala 71:55]
  wire  rsel_10 = _rsel_T[10]; // @[UserYanker.scala 71:55]
  wire  rsel_11 = _rsel_T[11]; // @[UserYanker.scala 71:55]
  wire  rsel_12 = _rsel_T[12]; // @[UserYanker.scala 71:55]
  wire  rsel_13 = _rsel_T[13]; // @[UserYanker.scala 71:55]
  wire  rsel_14 = _rsel_T[14]; // @[UserYanker.scala 71:55]
  wire  rsel_15 = _rsel_T[15]; // @[UserYanker.scala 71:55]
  wire  rsel_16 = _rsel_T[16]; // @[UserYanker.scala 71:55]
  wire  rsel_17 = _rsel_T[17]; // @[UserYanker.scala 71:55]
  wire  rsel_18 = _rsel_T[18]; // @[UserYanker.scala 71:55]
  wire  rsel_19 = _rsel_T[19]; // @[UserYanker.scala 71:55]
  wire  rsel_20 = _rsel_T[20]; // @[UserYanker.scala 71:55]
  wire  rsel_21 = _rsel_T[21]; // @[UserYanker.scala 71:55]
  wire  rsel_22 = _rsel_T[22]; // @[UserYanker.scala 71:55]
  wire  rsel_23 = _rsel_T[23]; // @[UserYanker.scala 71:55]
  wire  rsel_24 = _rsel_T[24]; // @[UserYanker.scala 71:55]
  wire  rsel_25 = _rsel_T[25]; // @[UserYanker.scala 71:55]
  wire  rsel_26 = _rsel_T[26]; // @[UserYanker.scala 71:55]
  wire  rsel_27 = _rsel_T[27]; // @[UserYanker.scala 71:55]
  wire  rsel_28 = _rsel_T[28]; // @[UserYanker.scala 71:55]
  wire  rsel_29 = _rsel_T[29]; // @[UserYanker.scala 71:55]
  wire  rsel_30 = _rsel_T[30]; // @[UserYanker.scala 71:55]
  wire  rsel_31 = _rsel_T[31]; // @[UserYanker.scala 71:55]
  wire  rsel_32 = _rsel_T[32]; // @[UserYanker.scala 71:55]
  wire  rsel_33 = _rsel_T[33]; // @[UserYanker.scala 71:55]
  wire  rsel_34 = _rsel_T[34]; // @[UserYanker.scala 71:55]
  wire  rsel_35 = _rsel_T[35]; // @[UserYanker.scala 71:55]
  wire  rsel_36 = _rsel_T[36]; // @[UserYanker.scala 71:55]
  wire  rsel_37 = _rsel_T[37]; // @[UserYanker.scala 71:55]
  wire  rsel_38 = _rsel_T[38]; // @[UserYanker.scala 71:55]
  wire  rsel_39 = _rsel_T[39]; // @[UserYanker.scala 71:55]
  wire  rsel_40 = _rsel_T[40]; // @[UserYanker.scala 71:55]
  wire  rsel_41 = _rsel_T[41]; // @[UserYanker.scala 71:55]
  wire  rsel_42 = _rsel_T[42]; // @[UserYanker.scala 71:55]
  wire  rsel_43 = _rsel_T[43]; // @[UserYanker.scala 71:55]
  wire  rsel_44 = _rsel_T[44]; // @[UserYanker.scala 71:55]
  wire  rsel_45 = _rsel_T[45]; // @[UserYanker.scala 71:55]
  wire  rsel_46 = _rsel_T[46]; // @[UserYanker.scala 71:55]
  wire  rsel_47 = _rsel_T[47]; // @[UserYanker.scala 71:55]
  wire  rsel_48 = _rsel_T[48]; // @[UserYanker.scala 71:55]
  wire  rsel_49 = _rsel_T[49]; // @[UserYanker.scala 71:55]
  wire  rsel_50 = _rsel_T[50]; // @[UserYanker.scala 71:55]
  wire  rsel_51 = _rsel_T[51]; // @[UserYanker.scala 71:55]
  wire  rsel_52 = _rsel_T[52]; // @[UserYanker.scala 71:55]
  wire  rsel_53 = _rsel_T[53]; // @[UserYanker.scala 71:55]
  wire  rsel_54 = _rsel_T[54]; // @[UserYanker.scala 71:55]
  wire  rsel_55 = _rsel_T[55]; // @[UserYanker.scala 71:55]
  wire  rsel_56 = _rsel_T[56]; // @[UserYanker.scala 71:55]
  wire  rsel_57 = _rsel_T[57]; // @[UserYanker.scala 71:55]
  wire  rsel_58 = _rsel_T[58]; // @[UserYanker.scala 71:55]
  wire  rsel_59 = _rsel_T[59]; // @[UserYanker.scala 71:55]
  wire  rsel_60 = _rsel_T[60]; // @[UserYanker.scala 71:55]
  wire  rsel_61 = _rsel_T[61]; // @[UserYanker.scala 71:55]
  wire  rsel_62 = _rsel_T[62]; // @[UserYanker.scala 71:55]
  wire  rsel_63 = _rsel_T[63]; // @[UserYanker.scala 71:55]
  wire  _aw_ready_WIRE_0 = Queue_64_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _aw_ready_WIRE_1 = Queue_65_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_321 = 6'h1 == auto_in_aw_bits_id ? _aw_ready_WIRE_1 : _aw_ready_WIRE_0; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_2 = Queue_66_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_322 = 6'h2 == auto_in_aw_bits_id ? _aw_ready_WIRE_2 : _GEN_321; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_3 = Queue_67_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_323 = 6'h3 == auto_in_aw_bits_id ? _aw_ready_WIRE_3 : _GEN_322; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_4 = Queue_68_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_324 = 6'h4 == auto_in_aw_bits_id ? _aw_ready_WIRE_4 : _GEN_323; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_5 = Queue_69_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_325 = 6'h5 == auto_in_aw_bits_id ? _aw_ready_WIRE_5 : _GEN_324; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_6 = Queue_70_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_326 = 6'h6 == auto_in_aw_bits_id ? _aw_ready_WIRE_6 : _GEN_325; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_7 = Queue_71_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_327 = 6'h7 == auto_in_aw_bits_id ? _aw_ready_WIRE_7 : _GEN_326; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_8 = Queue_72_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_328 = 6'h8 == auto_in_aw_bits_id ? _aw_ready_WIRE_8 : _GEN_327; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_9 = Queue_73_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_329 = 6'h9 == auto_in_aw_bits_id ? _aw_ready_WIRE_9 : _GEN_328; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_10 = Queue_74_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_330 = 6'ha == auto_in_aw_bits_id ? _aw_ready_WIRE_10 : _GEN_329; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_11 = Queue_75_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_331 = 6'hb == auto_in_aw_bits_id ? _aw_ready_WIRE_11 : _GEN_330; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_12 = Queue_76_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_332 = 6'hc == auto_in_aw_bits_id ? _aw_ready_WIRE_12 : _GEN_331; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_13 = Queue_77_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_333 = 6'hd == auto_in_aw_bits_id ? _aw_ready_WIRE_13 : _GEN_332; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_14 = Queue_78_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_334 = 6'he == auto_in_aw_bits_id ? _aw_ready_WIRE_14 : _GEN_333; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_15 = Queue_79_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_335 = 6'hf == auto_in_aw_bits_id ? _aw_ready_WIRE_15 : _GEN_334; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_16 = Queue_80_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_336 = 6'h10 == auto_in_aw_bits_id ? _aw_ready_WIRE_16 : _GEN_335; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_17 = Queue_81_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_337 = 6'h11 == auto_in_aw_bits_id ? _aw_ready_WIRE_17 : _GEN_336; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_18 = Queue_82_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_338 = 6'h12 == auto_in_aw_bits_id ? _aw_ready_WIRE_18 : _GEN_337; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_19 = Queue_83_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_339 = 6'h13 == auto_in_aw_bits_id ? _aw_ready_WIRE_19 : _GEN_338; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_20 = Queue_84_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_340 = 6'h14 == auto_in_aw_bits_id ? _aw_ready_WIRE_20 : _GEN_339; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_21 = Queue_85_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_341 = 6'h15 == auto_in_aw_bits_id ? _aw_ready_WIRE_21 : _GEN_340; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_22 = Queue_86_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_342 = 6'h16 == auto_in_aw_bits_id ? _aw_ready_WIRE_22 : _GEN_341; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_23 = Queue_87_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_343 = 6'h17 == auto_in_aw_bits_id ? _aw_ready_WIRE_23 : _GEN_342; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_24 = Queue_88_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_344 = 6'h18 == auto_in_aw_bits_id ? _aw_ready_WIRE_24 : _GEN_343; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_25 = Queue_89_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_345 = 6'h19 == auto_in_aw_bits_id ? _aw_ready_WIRE_25 : _GEN_344; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_26 = Queue_90_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_346 = 6'h1a == auto_in_aw_bits_id ? _aw_ready_WIRE_26 : _GEN_345; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_27 = Queue_91_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_347 = 6'h1b == auto_in_aw_bits_id ? _aw_ready_WIRE_27 : _GEN_346; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_28 = Queue_92_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_348 = 6'h1c == auto_in_aw_bits_id ? _aw_ready_WIRE_28 : _GEN_347; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_29 = Queue_93_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_349 = 6'h1d == auto_in_aw_bits_id ? _aw_ready_WIRE_29 : _GEN_348; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_30 = Queue_94_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_350 = 6'h1e == auto_in_aw_bits_id ? _aw_ready_WIRE_30 : _GEN_349; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_31 = Queue_95_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_351 = 6'h1f == auto_in_aw_bits_id ? _aw_ready_WIRE_31 : _GEN_350; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_32 = Queue_96_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_352 = 6'h20 == auto_in_aw_bits_id ? _aw_ready_WIRE_32 : _GEN_351; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_33 = Queue_97_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_353 = 6'h21 == auto_in_aw_bits_id ? _aw_ready_WIRE_33 : _GEN_352; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_34 = Queue_98_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_354 = 6'h22 == auto_in_aw_bits_id ? _aw_ready_WIRE_34 : _GEN_353; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_35 = Queue_99_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_355 = 6'h23 == auto_in_aw_bits_id ? _aw_ready_WIRE_35 : _GEN_354; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_36 = Queue_100_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_356 = 6'h24 == auto_in_aw_bits_id ? _aw_ready_WIRE_36 : _GEN_355; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_37 = Queue_101_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_357 = 6'h25 == auto_in_aw_bits_id ? _aw_ready_WIRE_37 : _GEN_356; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_38 = Queue_102_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_358 = 6'h26 == auto_in_aw_bits_id ? _aw_ready_WIRE_38 : _GEN_357; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_39 = Queue_103_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_359 = 6'h27 == auto_in_aw_bits_id ? _aw_ready_WIRE_39 : _GEN_358; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_40 = Queue_104_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_360 = 6'h28 == auto_in_aw_bits_id ? _aw_ready_WIRE_40 : _GEN_359; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_41 = Queue_105_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_361 = 6'h29 == auto_in_aw_bits_id ? _aw_ready_WIRE_41 : _GEN_360; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_42 = Queue_106_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_362 = 6'h2a == auto_in_aw_bits_id ? _aw_ready_WIRE_42 : _GEN_361; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_43 = Queue_107_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_363 = 6'h2b == auto_in_aw_bits_id ? _aw_ready_WIRE_43 : _GEN_362; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_44 = Queue_108_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_364 = 6'h2c == auto_in_aw_bits_id ? _aw_ready_WIRE_44 : _GEN_363; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_45 = Queue_109_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_365 = 6'h2d == auto_in_aw_bits_id ? _aw_ready_WIRE_45 : _GEN_364; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_46 = Queue_110_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_366 = 6'h2e == auto_in_aw_bits_id ? _aw_ready_WIRE_46 : _GEN_365; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_47 = Queue_111_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_367 = 6'h2f == auto_in_aw_bits_id ? _aw_ready_WIRE_47 : _GEN_366; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_48 = Queue_112_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_368 = 6'h30 == auto_in_aw_bits_id ? _aw_ready_WIRE_48 : _GEN_367; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_49 = Queue_113_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_369 = 6'h31 == auto_in_aw_bits_id ? _aw_ready_WIRE_49 : _GEN_368; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_50 = Queue_114_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_370 = 6'h32 == auto_in_aw_bits_id ? _aw_ready_WIRE_50 : _GEN_369; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_51 = Queue_115_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_371 = 6'h33 == auto_in_aw_bits_id ? _aw_ready_WIRE_51 : _GEN_370; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_52 = Queue_116_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_372 = 6'h34 == auto_in_aw_bits_id ? _aw_ready_WIRE_52 : _GEN_371; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_53 = Queue_117_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_373 = 6'h35 == auto_in_aw_bits_id ? _aw_ready_WIRE_53 : _GEN_372; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_54 = Queue_118_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_374 = 6'h36 == auto_in_aw_bits_id ? _aw_ready_WIRE_54 : _GEN_373; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_55 = Queue_119_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_375 = 6'h37 == auto_in_aw_bits_id ? _aw_ready_WIRE_55 : _GEN_374; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_56 = Queue_120_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_376 = 6'h38 == auto_in_aw_bits_id ? _aw_ready_WIRE_56 : _GEN_375; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_57 = Queue_121_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_377 = 6'h39 == auto_in_aw_bits_id ? _aw_ready_WIRE_57 : _GEN_376; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_58 = Queue_122_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_378 = 6'h3a == auto_in_aw_bits_id ? _aw_ready_WIRE_58 : _GEN_377; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_59 = Queue_123_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_379 = 6'h3b == auto_in_aw_bits_id ? _aw_ready_WIRE_59 : _GEN_378; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_60 = Queue_124_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_380 = 6'h3c == auto_in_aw_bits_id ? _aw_ready_WIRE_60 : _GEN_379; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_61 = Queue_125_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_381 = 6'h3d == auto_in_aw_bits_id ? _aw_ready_WIRE_61 : _GEN_380; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_62 = Queue_126_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_382 = 6'h3e == auto_in_aw_bits_id ? _aw_ready_WIRE_62 : _GEN_381; // @[UserYanker.scala 80:{36,36}]
  wire  _aw_ready_WIRE_63 = Queue_127_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_383 = 6'h3f == auto_in_aw_bits_id ? _aw_ready_WIRE_63 : _GEN_382; // @[UserYanker.scala 80:{36,36}]
  wire  _b_valid_WIRE_0 = Queue_64_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _b_valid_WIRE_1 = Queue_65_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_385 = 6'h1 == auto_out_b_bits_id ? _b_valid_WIRE_1 : _b_valid_WIRE_0; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_2 = Queue_66_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_386 = 6'h2 == auto_out_b_bits_id ? _b_valid_WIRE_2 : _GEN_385; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_3 = Queue_67_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_387 = 6'h3 == auto_out_b_bits_id ? _b_valid_WIRE_3 : _GEN_386; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_4 = Queue_68_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_388 = 6'h4 == auto_out_b_bits_id ? _b_valid_WIRE_4 : _GEN_387; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_5 = Queue_69_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_389 = 6'h5 == auto_out_b_bits_id ? _b_valid_WIRE_5 : _GEN_388; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_6 = Queue_70_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_390 = 6'h6 == auto_out_b_bits_id ? _b_valid_WIRE_6 : _GEN_389; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_7 = Queue_71_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_391 = 6'h7 == auto_out_b_bits_id ? _b_valid_WIRE_7 : _GEN_390; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_8 = Queue_72_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_392 = 6'h8 == auto_out_b_bits_id ? _b_valid_WIRE_8 : _GEN_391; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_9 = Queue_73_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_393 = 6'h9 == auto_out_b_bits_id ? _b_valid_WIRE_9 : _GEN_392; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_10 = Queue_74_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_394 = 6'ha == auto_out_b_bits_id ? _b_valid_WIRE_10 : _GEN_393; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_11 = Queue_75_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_395 = 6'hb == auto_out_b_bits_id ? _b_valid_WIRE_11 : _GEN_394; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_12 = Queue_76_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_396 = 6'hc == auto_out_b_bits_id ? _b_valid_WIRE_12 : _GEN_395; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_13 = Queue_77_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_397 = 6'hd == auto_out_b_bits_id ? _b_valid_WIRE_13 : _GEN_396; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_14 = Queue_78_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_398 = 6'he == auto_out_b_bits_id ? _b_valid_WIRE_14 : _GEN_397; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_15 = Queue_79_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_399 = 6'hf == auto_out_b_bits_id ? _b_valid_WIRE_15 : _GEN_398; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_16 = Queue_80_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_400 = 6'h10 == auto_out_b_bits_id ? _b_valid_WIRE_16 : _GEN_399; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_17 = Queue_81_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_401 = 6'h11 == auto_out_b_bits_id ? _b_valid_WIRE_17 : _GEN_400; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_18 = Queue_82_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_402 = 6'h12 == auto_out_b_bits_id ? _b_valid_WIRE_18 : _GEN_401; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_19 = Queue_83_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_403 = 6'h13 == auto_out_b_bits_id ? _b_valid_WIRE_19 : _GEN_402; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_20 = Queue_84_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_404 = 6'h14 == auto_out_b_bits_id ? _b_valid_WIRE_20 : _GEN_403; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_21 = Queue_85_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_405 = 6'h15 == auto_out_b_bits_id ? _b_valid_WIRE_21 : _GEN_404; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_22 = Queue_86_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_406 = 6'h16 == auto_out_b_bits_id ? _b_valid_WIRE_22 : _GEN_405; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_23 = Queue_87_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_407 = 6'h17 == auto_out_b_bits_id ? _b_valid_WIRE_23 : _GEN_406; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_24 = Queue_88_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_408 = 6'h18 == auto_out_b_bits_id ? _b_valid_WIRE_24 : _GEN_407; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_25 = Queue_89_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_409 = 6'h19 == auto_out_b_bits_id ? _b_valid_WIRE_25 : _GEN_408; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_26 = Queue_90_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_410 = 6'h1a == auto_out_b_bits_id ? _b_valid_WIRE_26 : _GEN_409; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_27 = Queue_91_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_411 = 6'h1b == auto_out_b_bits_id ? _b_valid_WIRE_27 : _GEN_410; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_28 = Queue_92_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_412 = 6'h1c == auto_out_b_bits_id ? _b_valid_WIRE_28 : _GEN_411; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_29 = Queue_93_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_413 = 6'h1d == auto_out_b_bits_id ? _b_valid_WIRE_29 : _GEN_412; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_30 = Queue_94_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_414 = 6'h1e == auto_out_b_bits_id ? _b_valid_WIRE_30 : _GEN_413; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_31 = Queue_95_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_415 = 6'h1f == auto_out_b_bits_id ? _b_valid_WIRE_31 : _GEN_414; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_32 = Queue_96_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_416 = 6'h20 == auto_out_b_bits_id ? _b_valid_WIRE_32 : _GEN_415; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_33 = Queue_97_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_417 = 6'h21 == auto_out_b_bits_id ? _b_valid_WIRE_33 : _GEN_416; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_34 = Queue_98_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_418 = 6'h22 == auto_out_b_bits_id ? _b_valid_WIRE_34 : _GEN_417; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_35 = Queue_99_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_419 = 6'h23 == auto_out_b_bits_id ? _b_valid_WIRE_35 : _GEN_418; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_36 = Queue_100_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_420 = 6'h24 == auto_out_b_bits_id ? _b_valid_WIRE_36 : _GEN_419; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_37 = Queue_101_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_421 = 6'h25 == auto_out_b_bits_id ? _b_valid_WIRE_37 : _GEN_420; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_38 = Queue_102_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_422 = 6'h26 == auto_out_b_bits_id ? _b_valid_WIRE_38 : _GEN_421; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_39 = Queue_103_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_423 = 6'h27 == auto_out_b_bits_id ? _b_valid_WIRE_39 : _GEN_422; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_40 = Queue_104_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_424 = 6'h28 == auto_out_b_bits_id ? _b_valid_WIRE_40 : _GEN_423; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_41 = Queue_105_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_425 = 6'h29 == auto_out_b_bits_id ? _b_valid_WIRE_41 : _GEN_424; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_42 = Queue_106_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_426 = 6'h2a == auto_out_b_bits_id ? _b_valid_WIRE_42 : _GEN_425; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_43 = Queue_107_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_427 = 6'h2b == auto_out_b_bits_id ? _b_valid_WIRE_43 : _GEN_426; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_44 = Queue_108_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_428 = 6'h2c == auto_out_b_bits_id ? _b_valid_WIRE_44 : _GEN_427; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_45 = Queue_109_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_429 = 6'h2d == auto_out_b_bits_id ? _b_valid_WIRE_45 : _GEN_428; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_46 = Queue_110_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_430 = 6'h2e == auto_out_b_bits_id ? _b_valid_WIRE_46 : _GEN_429; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_47 = Queue_111_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_431 = 6'h2f == auto_out_b_bits_id ? _b_valid_WIRE_47 : _GEN_430; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_48 = Queue_112_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_432 = 6'h30 == auto_out_b_bits_id ? _b_valid_WIRE_48 : _GEN_431; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_49 = Queue_113_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_433 = 6'h31 == auto_out_b_bits_id ? _b_valid_WIRE_49 : _GEN_432; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_50 = Queue_114_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_434 = 6'h32 == auto_out_b_bits_id ? _b_valid_WIRE_50 : _GEN_433; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_51 = Queue_115_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_435 = 6'h33 == auto_out_b_bits_id ? _b_valid_WIRE_51 : _GEN_434; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_52 = Queue_116_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_436 = 6'h34 == auto_out_b_bits_id ? _b_valid_WIRE_52 : _GEN_435; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_53 = Queue_117_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_437 = 6'h35 == auto_out_b_bits_id ? _b_valid_WIRE_53 : _GEN_436; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_54 = Queue_118_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_438 = 6'h36 == auto_out_b_bits_id ? _b_valid_WIRE_54 : _GEN_437; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_55 = Queue_119_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_439 = 6'h37 == auto_out_b_bits_id ? _b_valid_WIRE_55 : _GEN_438; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_56 = Queue_120_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_440 = 6'h38 == auto_out_b_bits_id ? _b_valid_WIRE_56 : _GEN_439; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_57 = Queue_121_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_441 = 6'h39 == auto_out_b_bits_id ? _b_valid_WIRE_57 : _GEN_440; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_58 = Queue_122_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_442 = 6'h3a == auto_out_b_bits_id ? _b_valid_WIRE_58 : _GEN_441; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_59 = Queue_123_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_443 = 6'h3b == auto_out_b_bits_id ? _b_valid_WIRE_59 : _GEN_442; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_60 = Queue_124_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_444 = 6'h3c == auto_out_b_bits_id ? _b_valid_WIRE_60 : _GEN_443; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_61 = Queue_125_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_445 = 6'h3d == auto_out_b_bits_id ? _b_valid_WIRE_61 : _GEN_444; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_62 = Queue_126_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_446 = 6'h3e == auto_out_b_bits_id ? _b_valid_WIRE_62 : _GEN_445; // @[UserYanker.scala 87:{28,28}]
  wire  _b_valid_WIRE_63 = Queue_127_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_447 = 6'h3f == auto_out_b_bits_id ? _b_valid_WIRE_63 : _GEN_446; // @[UserYanker.scala 87:{28,28}]
  wire [1:0] _b_bits_WIRE_0_extra_id = Queue_64_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _b_bits_WIRE_1_extra_id = Queue_65_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_449 = 6'h1 == auto_out_b_bits_id ? _b_bits_WIRE_1_extra_id : _b_bits_WIRE_0_extra_id; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_2_extra_id = Queue_66_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_450 = 6'h2 == auto_out_b_bits_id ? _b_bits_WIRE_2_extra_id : _GEN_449; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_3_extra_id = Queue_67_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_451 = 6'h3 == auto_out_b_bits_id ? _b_bits_WIRE_3_extra_id : _GEN_450; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_4_extra_id = Queue_68_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_452 = 6'h4 == auto_out_b_bits_id ? _b_bits_WIRE_4_extra_id : _GEN_451; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_5_extra_id = Queue_69_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_453 = 6'h5 == auto_out_b_bits_id ? _b_bits_WIRE_5_extra_id : _GEN_452; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_6_extra_id = Queue_70_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_454 = 6'h6 == auto_out_b_bits_id ? _b_bits_WIRE_6_extra_id : _GEN_453; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_7_extra_id = Queue_71_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_455 = 6'h7 == auto_out_b_bits_id ? _b_bits_WIRE_7_extra_id : _GEN_454; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_8_extra_id = Queue_72_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_456 = 6'h8 == auto_out_b_bits_id ? _b_bits_WIRE_8_extra_id : _GEN_455; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_9_extra_id = Queue_73_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_457 = 6'h9 == auto_out_b_bits_id ? _b_bits_WIRE_9_extra_id : _GEN_456; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_10_extra_id = Queue_74_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_458 = 6'ha == auto_out_b_bits_id ? _b_bits_WIRE_10_extra_id : _GEN_457; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_11_extra_id = Queue_75_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_459 = 6'hb == auto_out_b_bits_id ? _b_bits_WIRE_11_extra_id : _GEN_458; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_12_extra_id = Queue_76_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_460 = 6'hc == auto_out_b_bits_id ? _b_bits_WIRE_12_extra_id : _GEN_459; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_13_extra_id = Queue_77_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_461 = 6'hd == auto_out_b_bits_id ? _b_bits_WIRE_13_extra_id : _GEN_460; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_14_extra_id = Queue_78_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_462 = 6'he == auto_out_b_bits_id ? _b_bits_WIRE_14_extra_id : _GEN_461; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_15_extra_id = Queue_79_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_463 = 6'hf == auto_out_b_bits_id ? _b_bits_WIRE_15_extra_id : _GEN_462; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_16_extra_id = Queue_80_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_464 = 6'h10 == auto_out_b_bits_id ? _b_bits_WIRE_16_extra_id : _GEN_463; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_17_extra_id = Queue_81_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_465 = 6'h11 == auto_out_b_bits_id ? _b_bits_WIRE_17_extra_id : _GEN_464; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_18_extra_id = Queue_82_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_466 = 6'h12 == auto_out_b_bits_id ? _b_bits_WIRE_18_extra_id : _GEN_465; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_19_extra_id = Queue_83_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_467 = 6'h13 == auto_out_b_bits_id ? _b_bits_WIRE_19_extra_id : _GEN_466; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_20_extra_id = Queue_84_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_468 = 6'h14 == auto_out_b_bits_id ? _b_bits_WIRE_20_extra_id : _GEN_467; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_21_extra_id = Queue_85_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_469 = 6'h15 == auto_out_b_bits_id ? _b_bits_WIRE_21_extra_id : _GEN_468; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_22_extra_id = Queue_86_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_470 = 6'h16 == auto_out_b_bits_id ? _b_bits_WIRE_22_extra_id : _GEN_469; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_23_extra_id = Queue_87_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_471 = 6'h17 == auto_out_b_bits_id ? _b_bits_WIRE_23_extra_id : _GEN_470; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_24_extra_id = Queue_88_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_472 = 6'h18 == auto_out_b_bits_id ? _b_bits_WIRE_24_extra_id : _GEN_471; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_25_extra_id = Queue_89_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_473 = 6'h19 == auto_out_b_bits_id ? _b_bits_WIRE_25_extra_id : _GEN_472; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_26_extra_id = Queue_90_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_474 = 6'h1a == auto_out_b_bits_id ? _b_bits_WIRE_26_extra_id : _GEN_473; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_27_extra_id = Queue_91_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_475 = 6'h1b == auto_out_b_bits_id ? _b_bits_WIRE_27_extra_id : _GEN_474; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_28_extra_id = Queue_92_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_476 = 6'h1c == auto_out_b_bits_id ? _b_bits_WIRE_28_extra_id : _GEN_475; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_29_extra_id = Queue_93_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_477 = 6'h1d == auto_out_b_bits_id ? _b_bits_WIRE_29_extra_id : _GEN_476; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_30_extra_id = Queue_94_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_478 = 6'h1e == auto_out_b_bits_id ? _b_bits_WIRE_30_extra_id : _GEN_477; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_31_extra_id = Queue_95_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_479 = 6'h1f == auto_out_b_bits_id ? _b_bits_WIRE_31_extra_id : _GEN_478; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_32_extra_id = Queue_96_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_480 = 6'h20 == auto_out_b_bits_id ? _b_bits_WIRE_32_extra_id : _GEN_479; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_33_extra_id = Queue_97_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_481 = 6'h21 == auto_out_b_bits_id ? _b_bits_WIRE_33_extra_id : _GEN_480; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_34_extra_id = Queue_98_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_482 = 6'h22 == auto_out_b_bits_id ? _b_bits_WIRE_34_extra_id : _GEN_481; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_35_extra_id = Queue_99_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_483 = 6'h23 == auto_out_b_bits_id ? _b_bits_WIRE_35_extra_id : _GEN_482; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_36_extra_id = Queue_100_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_484 = 6'h24 == auto_out_b_bits_id ? _b_bits_WIRE_36_extra_id : _GEN_483; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_37_extra_id = Queue_101_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_485 = 6'h25 == auto_out_b_bits_id ? _b_bits_WIRE_37_extra_id : _GEN_484; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_38_extra_id = Queue_102_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_486 = 6'h26 == auto_out_b_bits_id ? _b_bits_WIRE_38_extra_id : _GEN_485; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_39_extra_id = Queue_103_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_487 = 6'h27 == auto_out_b_bits_id ? _b_bits_WIRE_39_extra_id : _GEN_486; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_40_extra_id = Queue_104_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_488 = 6'h28 == auto_out_b_bits_id ? _b_bits_WIRE_40_extra_id : _GEN_487; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_41_extra_id = Queue_105_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_489 = 6'h29 == auto_out_b_bits_id ? _b_bits_WIRE_41_extra_id : _GEN_488; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_42_extra_id = Queue_106_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_490 = 6'h2a == auto_out_b_bits_id ? _b_bits_WIRE_42_extra_id : _GEN_489; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_43_extra_id = Queue_107_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_491 = 6'h2b == auto_out_b_bits_id ? _b_bits_WIRE_43_extra_id : _GEN_490; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_44_extra_id = Queue_108_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_492 = 6'h2c == auto_out_b_bits_id ? _b_bits_WIRE_44_extra_id : _GEN_491; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_45_extra_id = Queue_109_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_493 = 6'h2d == auto_out_b_bits_id ? _b_bits_WIRE_45_extra_id : _GEN_492; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_46_extra_id = Queue_110_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_494 = 6'h2e == auto_out_b_bits_id ? _b_bits_WIRE_46_extra_id : _GEN_493; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_47_extra_id = Queue_111_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_495 = 6'h2f == auto_out_b_bits_id ? _b_bits_WIRE_47_extra_id : _GEN_494; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_48_extra_id = Queue_112_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_496 = 6'h30 == auto_out_b_bits_id ? _b_bits_WIRE_48_extra_id : _GEN_495; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_49_extra_id = Queue_113_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_497 = 6'h31 == auto_out_b_bits_id ? _b_bits_WIRE_49_extra_id : _GEN_496; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_50_extra_id = Queue_114_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_498 = 6'h32 == auto_out_b_bits_id ? _b_bits_WIRE_50_extra_id : _GEN_497; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_51_extra_id = Queue_115_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_499 = 6'h33 == auto_out_b_bits_id ? _b_bits_WIRE_51_extra_id : _GEN_498; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_52_extra_id = Queue_116_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_500 = 6'h34 == auto_out_b_bits_id ? _b_bits_WIRE_52_extra_id : _GEN_499; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_53_extra_id = Queue_117_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_501 = 6'h35 == auto_out_b_bits_id ? _b_bits_WIRE_53_extra_id : _GEN_500; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_54_extra_id = Queue_118_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_502 = 6'h36 == auto_out_b_bits_id ? _b_bits_WIRE_54_extra_id : _GEN_501; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_55_extra_id = Queue_119_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_503 = 6'h37 == auto_out_b_bits_id ? _b_bits_WIRE_55_extra_id : _GEN_502; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_56_extra_id = Queue_120_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_504 = 6'h38 == auto_out_b_bits_id ? _b_bits_WIRE_56_extra_id : _GEN_503; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_57_extra_id = Queue_121_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_505 = 6'h39 == auto_out_b_bits_id ? _b_bits_WIRE_57_extra_id : _GEN_504; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_58_extra_id = Queue_122_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_506 = 6'h3a == auto_out_b_bits_id ? _b_bits_WIRE_58_extra_id : _GEN_505; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_59_extra_id = Queue_123_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_507 = 6'h3b == auto_out_b_bits_id ? _b_bits_WIRE_59_extra_id : _GEN_506; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_60_extra_id = Queue_124_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_508 = 6'h3c == auto_out_b_bits_id ? _b_bits_WIRE_60_extra_id : _GEN_507; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_61_extra_id = Queue_125_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_509 = 6'h3d == auto_out_b_bits_id ? _b_bits_WIRE_61_extra_id : _GEN_508; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_62_extra_id = Queue_126_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _GEN_510 = 6'h3e == auto_out_b_bits_id ? _b_bits_WIRE_62_extra_id : _GEN_509; // @[BundleMap.scala 247:{19,19}]
  wire [1:0] _b_bits_WIRE_63_extra_id = Queue_127_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _b_bits_WIRE_0_tl_state_source = Queue_64_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _b_bits_WIRE_1_tl_state_source = Queue_65_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_513 = 6'h1 == auto_out_b_bits_id ? _b_bits_WIRE_1_tl_state_source : _b_bits_WIRE_0_tl_state_source; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_2_tl_state_source = Queue_66_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_514 = 6'h2 == auto_out_b_bits_id ? _b_bits_WIRE_2_tl_state_source : _GEN_513; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_3_tl_state_source = Queue_67_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_515 = 6'h3 == auto_out_b_bits_id ? _b_bits_WIRE_3_tl_state_source : _GEN_514; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_4_tl_state_source = Queue_68_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_516 = 6'h4 == auto_out_b_bits_id ? _b_bits_WIRE_4_tl_state_source : _GEN_515; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_5_tl_state_source = Queue_69_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_517 = 6'h5 == auto_out_b_bits_id ? _b_bits_WIRE_5_tl_state_source : _GEN_516; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_6_tl_state_source = Queue_70_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_518 = 6'h6 == auto_out_b_bits_id ? _b_bits_WIRE_6_tl_state_source : _GEN_517; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_7_tl_state_source = Queue_71_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_519 = 6'h7 == auto_out_b_bits_id ? _b_bits_WIRE_7_tl_state_source : _GEN_518; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_8_tl_state_source = Queue_72_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_520 = 6'h8 == auto_out_b_bits_id ? _b_bits_WIRE_8_tl_state_source : _GEN_519; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_9_tl_state_source = Queue_73_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_521 = 6'h9 == auto_out_b_bits_id ? _b_bits_WIRE_9_tl_state_source : _GEN_520; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_10_tl_state_source = Queue_74_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_522 = 6'ha == auto_out_b_bits_id ? _b_bits_WIRE_10_tl_state_source : _GEN_521; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_11_tl_state_source = Queue_75_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_523 = 6'hb == auto_out_b_bits_id ? _b_bits_WIRE_11_tl_state_source : _GEN_522; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_12_tl_state_source = Queue_76_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_524 = 6'hc == auto_out_b_bits_id ? _b_bits_WIRE_12_tl_state_source : _GEN_523; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_13_tl_state_source = Queue_77_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_525 = 6'hd == auto_out_b_bits_id ? _b_bits_WIRE_13_tl_state_source : _GEN_524; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_14_tl_state_source = Queue_78_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_526 = 6'he == auto_out_b_bits_id ? _b_bits_WIRE_14_tl_state_source : _GEN_525; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_15_tl_state_source = Queue_79_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_527 = 6'hf == auto_out_b_bits_id ? _b_bits_WIRE_15_tl_state_source : _GEN_526; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_16_tl_state_source = Queue_80_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_528 = 6'h10 == auto_out_b_bits_id ? _b_bits_WIRE_16_tl_state_source : _GEN_527; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_17_tl_state_source = Queue_81_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_529 = 6'h11 == auto_out_b_bits_id ? _b_bits_WIRE_17_tl_state_source : _GEN_528; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_18_tl_state_source = Queue_82_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_530 = 6'h12 == auto_out_b_bits_id ? _b_bits_WIRE_18_tl_state_source : _GEN_529; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_19_tl_state_source = Queue_83_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_531 = 6'h13 == auto_out_b_bits_id ? _b_bits_WIRE_19_tl_state_source : _GEN_530; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_20_tl_state_source = Queue_84_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_532 = 6'h14 == auto_out_b_bits_id ? _b_bits_WIRE_20_tl_state_source : _GEN_531; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_21_tl_state_source = Queue_85_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_533 = 6'h15 == auto_out_b_bits_id ? _b_bits_WIRE_21_tl_state_source : _GEN_532; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_22_tl_state_source = Queue_86_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_534 = 6'h16 == auto_out_b_bits_id ? _b_bits_WIRE_22_tl_state_source : _GEN_533; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_23_tl_state_source = Queue_87_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_535 = 6'h17 == auto_out_b_bits_id ? _b_bits_WIRE_23_tl_state_source : _GEN_534; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_24_tl_state_source = Queue_88_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_536 = 6'h18 == auto_out_b_bits_id ? _b_bits_WIRE_24_tl_state_source : _GEN_535; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_25_tl_state_source = Queue_89_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_537 = 6'h19 == auto_out_b_bits_id ? _b_bits_WIRE_25_tl_state_source : _GEN_536; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_26_tl_state_source = Queue_90_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_538 = 6'h1a == auto_out_b_bits_id ? _b_bits_WIRE_26_tl_state_source : _GEN_537; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_27_tl_state_source = Queue_91_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_539 = 6'h1b == auto_out_b_bits_id ? _b_bits_WIRE_27_tl_state_source : _GEN_538; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_28_tl_state_source = Queue_92_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_540 = 6'h1c == auto_out_b_bits_id ? _b_bits_WIRE_28_tl_state_source : _GEN_539; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_29_tl_state_source = Queue_93_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_541 = 6'h1d == auto_out_b_bits_id ? _b_bits_WIRE_29_tl_state_source : _GEN_540; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_30_tl_state_source = Queue_94_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_542 = 6'h1e == auto_out_b_bits_id ? _b_bits_WIRE_30_tl_state_source : _GEN_541; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_31_tl_state_source = Queue_95_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_543 = 6'h1f == auto_out_b_bits_id ? _b_bits_WIRE_31_tl_state_source : _GEN_542; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_32_tl_state_source = Queue_96_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_544 = 6'h20 == auto_out_b_bits_id ? _b_bits_WIRE_32_tl_state_source : _GEN_543; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_33_tl_state_source = Queue_97_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_545 = 6'h21 == auto_out_b_bits_id ? _b_bits_WIRE_33_tl_state_source : _GEN_544; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_34_tl_state_source = Queue_98_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_546 = 6'h22 == auto_out_b_bits_id ? _b_bits_WIRE_34_tl_state_source : _GEN_545; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_35_tl_state_source = Queue_99_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_547 = 6'h23 == auto_out_b_bits_id ? _b_bits_WIRE_35_tl_state_source : _GEN_546; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_36_tl_state_source = Queue_100_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_548 = 6'h24 == auto_out_b_bits_id ? _b_bits_WIRE_36_tl_state_source : _GEN_547; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_37_tl_state_source = Queue_101_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_549 = 6'h25 == auto_out_b_bits_id ? _b_bits_WIRE_37_tl_state_source : _GEN_548; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_38_tl_state_source = Queue_102_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_550 = 6'h26 == auto_out_b_bits_id ? _b_bits_WIRE_38_tl_state_source : _GEN_549; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_39_tl_state_source = Queue_103_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_551 = 6'h27 == auto_out_b_bits_id ? _b_bits_WIRE_39_tl_state_source : _GEN_550; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_40_tl_state_source = Queue_104_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_552 = 6'h28 == auto_out_b_bits_id ? _b_bits_WIRE_40_tl_state_source : _GEN_551; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_41_tl_state_source = Queue_105_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_553 = 6'h29 == auto_out_b_bits_id ? _b_bits_WIRE_41_tl_state_source : _GEN_552; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_42_tl_state_source = Queue_106_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_554 = 6'h2a == auto_out_b_bits_id ? _b_bits_WIRE_42_tl_state_source : _GEN_553; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_43_tl_state_source = Queue_107_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_555 = 6'h2b == auto_out_b_bits_id ? _b_bits_WIRE_43_tl_state_source : _GEN_554; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_44_tl_state_source = Queue_108_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_556 = 6'h2c == auto_out_b_bits_id ? _b_bits_WIRE_44_tl_state_source : _GEN_555; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_45_tl_state_source = Queue_109_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_557 = 6'h2d == auto_out_b_bits_id ? _b_bits_WIRE_45_tl_state_source : _GEN_556; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_46_tl_state_source = Queue_110_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_558 = 6'h2e == auto_out_b_bits_id ? _b_bits_WIRE_46_tl_state_source : _GEN_557; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_47_tl_state_source = Queue_111_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_559 = 6'h2f == auto_out_b_bits_id ? _b_bits_WIRE_47_tl_state_source : _GEN_558; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_48_tl_state_source = Queue_112_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_560 = 6'h30 == auto_out_b_bits_id ? _b_bits_WIRE_48_tl_state_source : _GEN_559; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_49_tl_state_source = Queue_113_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_561 = 6'h31 == auto_out_b_bits_id ? _b_bits_WIRE_49_tl_state_source : _GEN_560; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_50_tl_state_source = Queue_114_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_562 = 6'h32 == auto_out_b_bits_id ? _b_bits_WIRE_50_tl_state_source : _GEN_561; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_51_tl_state_source = Queue_115_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_563 = 6'h33 == auto_out_b_bits_id ? _b_bits_WIRE_51_tl_state_source : _GEN_562; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_52_tl_state_source = Queue_116_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_564 = 6'h34 == auto_out_b_bits_id ? _b_bits_WIRE_52_tl_state_source : _GEN_563; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_53_tl_state_source = Queue_117_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_565 = 6'h35 == auto_out_b_bits_id ? _b_bits_WIRE_53_tl_state_source : _GEN_564; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_54_tl_state_source = Queue_118_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_566 = 6'h36 == auto_out_b_bits_id ? _b_bits_WIRE_54_tl_state_source : _GEN_565; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_55_tl_state_source = Queue_119_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_567 = 6'h37 == auto_out_b_bits_id ? _b_bits_WIRE_55_tl_state_source : _GEN_566; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_56_tl_state_source = Queue_120_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_568 = 6'h38 == auto_out_b_bits_id ? _b_bits_WIRE_56_tl_state_source : _GEN_567; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_57_tl_state_source = Queue_121_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_569 = 6'h39 == auto_out_b_bits_id ? _b_bits_WIRE_57_tl_state_source : _GEN_568; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_58_tl_state_source = Queue_122_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_570 = 6'h3a == auto_out_b_bits_id ? _b_bits_WIRE_58_tl_state_source : _GEN_569; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_59_tl_state_source = Queue_123_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_571 = 6'h3b == auto_out_b_bits_id ? _b_bits_WIRE_59_tl_state_source : _GEN_570; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_60_tl_state_source = Queue_124_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_572 = 6'h3c == auto_out_b_bits_id ? _b_bits_WIRE_60_tl_state_source : _GEN_571; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_61_tl_state_source = Queue_125_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_573 = 6'h3d == auto_out_b_bits_id ? _b_bits_WIRE_61_tl_state_source : _GEN_572; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_62_tl_state_source = Queue_126_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [6:0] _GEN_574 = 6'h3e == auto_out_b_bits_id ? _b_bits_WIRE_62_tl_state_source : _GEN_573; // @[BundleMap.scala 247:{19,19}]
  wire [6:0] _b_bits_WIRE_63_tl_state_source = Queue_127_io_deq_bits_tl_state_source; // @[UserYanker.scala 86:{27,27}]
  wire [63:0] _awsel_T = 64'h1 << auto_in_aw_bits_id; // @[OneHot.scala 64:12]
  wire  awsel_0 = _awsel_T[0]; // @[UserYanker.scala 91:55]
  wire  awsel_1 = _awsel_T[1]; // @[UserYanker.scala 91:55]
  wire  awsel_2 = _awsel_T[2]; // @[UserYanker.scala 91:55]
  wire  awsel_3 = _awsel_T[3]; // @[UserYanker.scala 91:55]
  wire  awsel_4 = _awsel_T[4]; // @[UserYanker.scala 91:55]
  wire  awsel_5 = _awsel_T[5]; // @[UserYanker.scala 91:55]
  wire  awsel_6 = _awsel_T[6]; // @[UserYanker.scala 91:55]
  wire  awsel_7 = _awsel_T[7]; // @[UserYanker.scala 91:55]
  wire  awsel_8 = _awsel_T[8]; // @[UserYanker.scala 91:55]
  wire  awsel_9 = _awsel_T[9]; // @[UserYanker.scala 91:55]
  wire  awsel_10 = _awsel_T[10]; // @[UserYanker.scala 91:55]
  wire  awsel_11 = _awsel_T[11]; // @[UserYanker.scala 91:55]
  wire  awsel_12 = _awsel_T[12]; // @[UserYanker.scala 91:55]
  wire  awsel_13 = _awsel_T[13]; // @[UserYanker.scala 91:55]
  wire  awsel_14 = _awsel_T[14]; // @[UserYanker.scala 91:55]
  wire  awsel_15 = _awsel_T[15]; // @[UserYanker.scala 91:55]
  wire  awsel_16 = _awsel_T[16]; // @[UserYanker.scala 91:55]
  wire  awsel_17 = _awsel_T[17]; // @[UserYanker.scala 91:55]
  wire  awsel_18 = _awsel_T[18]; // @[UserYanker.scala 91:55]
  wire  awsel_19 = _awsel_T[19]; // @[UserYanker.scala 91:55]
  wire  awsel_20 = _awsel_T[20]; // @[UserYanker.scala 91:55]
  wire  awsel_21 = _awsel_T[21]; // @[UserYanker.scala 91:55]
  wire  awsel_22 = _awsel_T[22]; // @[UserYanker.scala 91:55]
  wire  awsel_23 = _awsel_T[23]; // @[UserYanker.scala 91:55]
  wire  awsel_24 = _awsel_T[24]; // @[UserYanker.scala 91:55]
  wire  awsel_25 = _awsel_T[25]; // @[UserYanker.scala 91:55]
  wire  awsel_26 = _awsel_T[26]; // @[UserYanker.scala 91:55]
  wire  awsel_27 = _awsel_T[27]; // @[UserYanker.scala 91:55]
  wire  awsel_28 = _awsel_T[28]; // @[UserYanker.scala 91:55]
  wire  awsel_29 = _awsel_T[29]; // @[UserYanker.scala 91:55]
  wire  awsel_30 = _awsel_T[30]; // @[UserYanker.scala 91:55]
  wire  awsel_31 = _awsel_T[31]; // @[UserYanker.scala 91:55]
  wire  awsel_32 = _awsel_T[32]; // @[UserYanker.scala 91:55]
  wire  awsel_33 = _awsel_T[33]; // @[UserYanker.scala 91:55]
  wire  awsel_34 = _awsel_T[34]; // @[UserYanker.scala 91:55]
  wire  awsel_35 = _awsel_T[35]; // @[UserYanker.scala 91:55]
  wire  awsel_36 = _awsel_T[36]; // @[UserYanker.scala 91:55]
  wire  awsel_37 = _awsel_T[37]; // @[UserYanker.scala 91:55]
  wire  awsel_38 = _awsel_T[38]; // @[UserYanker.scala 91:55]
  wire  awsel_39 = _awsel_T[39]; // @[UserYanker.scala 91:55]
  wire  awsel_40 = _awsel_T[40]; // @[UserYanker.scala 91:55]
  wire  awsel_41 = _awsel_T[41]; // @[UserYanker.scala 91:55]
  wire  awsel_42 = _awsel_T[42]; // @[UserYanker.scala 91:55]
  wire  awsel_43 = _awsel_T[43]; // @[UserYanker.scala 91:55]
  wire  awsel_44 = _awsel_T[44]; // @[UserYanker.scala 91:55]
  wire  awsel_45 = _awsel_T[45]; // @[UserYanker.scala 91:55]
  wire  awsel_46 = _awsel_T[46]; // @[UserYanker.scala 91:55]
  wire  awsel_47 = _awsel_T[47]; // @[UserYanker.scala 91:55]
  wire  awsel_48 = _awsel_T[48]; // @[UserYanker.scala 91:55]
  wire  awsel_49 = _awsel_T[49]; // @[UserYanker.scala 91:55]
  wire  awsel_50 = _awsel_T[50]; // @[UserYanker.scala 91:55]
  wire  awsel_51 = _awsel_T[51]; // @[UserYanker.scala 91:55]
  wire  awsel_52 = _awsel_T[52]; // @[UserYanker.scala 91:55]
  wire  awsel_53 = _awsel_T[53]; // @[UserYanker.scala 91:55]
  wire  awsel_54 = _awsel_T[54]; // @[UserYanker.scala 91:55]
  wire  awsel_55 = _awsel_T[55]; // @[UserYanker.scala 91:55]
  wire  awsel_56 = _awsel_T[56]; // @[UserYanker.scala 91:55]
  wire  awsel_57 = _awsel_T[57]; // @[UserYanker.scala 91:55]
  wire  awsel_58 = _awsel_T[58]; // @[UserYanker.scala 91:55]
  wire  awsel_59 = _awsel_T[59]; // @[UserYanker.scala 91:55]
  wire  awsel_60 = _awsel_T[60]; // @[UserYanker.scala 91:55]
  wire  awsel_61 = _awsel_T[61]; // @[UserYanker.scala 91:55]
  wire  awsel_62 = _awsel_T[62]; // @[UserYanker.scala 91:55]
  wire  awsel_63 = _awsel_T[63]; // @[UserYanker.scala 91:55]
  wire [63:0] _bsel_T = 64'h1 << auto_out_b_bits_id; // @[OneHot.scala 64:12]
  wire  bsel_0 = _bsel_T[0]; // @[UserYanker.scala 92:55]
  wire  bsel_1 = _bsel_T[1]; // @[UserYanker.scala 92:55]
  wire  bsel_2 = _bsel_T[2]; // @[UserYanker.scala 92:55]
  wire  bsel_3 = _bsel_T[3]; // @[UserYanker.scala 92:55]
  wire  bsel_4 = _bsel_T[4]; // @[UserYanker.scala 92:55]
  wire  bsel_5 = _bsel_T[5]; // @[UserYanker.scala 92:55]
  wire  bsel_6 = _bsel_T[6]; // @[UserYanker.scala 92:55]
  wire  bsel_7 = _bsel_T[7]; // @[UserYanker.scala 92:55]
  wire  bsel_8 = _bsel_T[8]; // @[UserYanker.scala 92:55]
  wire  bsel_9 = _bsel_T[9]; // @[UserYanker.scala 92:55]
  wire  bsel_10 = _bsel_T[10]; // @[UserYanker.scala 92:55]
  wire  bsel_11 = _bsel_T[11]; // @[UserYanker.scala 92:55]
  wire  bsel_12 = _bsel_T[12]; // @[UserYanker.scala 92:55]
  wire  bsel_13 = _bsel_T[13]; // @[UserYanker.scala 92:55]
  wire  bsel_14 = _bsel_T[14]; // @[UserYanker.scala 92:55]
  wire  bsel_15 = _bsel_T[15]; // @[UserYanker.scala 92:55]
  wire  bsel_16 = _bsel_T[16]; // @[UserYanker.scala 92:55]
  wire  bsel_17 = _bsel_T[17]; // @[UserYanker.scala 92:55]
  wire  bsel_18 = _bsel_T[18]; // @[UserYanker.scala 92:55]
  wire  bsel_19 = _bsel_T[19]; // @[UserYanker.scala 92:55]
  wire  bsel_20 = _bsel_T[20]; // @[UserYanker.scala 92:55]
  wire  bsel_21 = _bsel_T[21]; // @[UserYanker.scala 92:55]
  wire  bsel_22 = _bsel_T[22]; // @[UserYanker.scala 92:55]
  wire  bsel_23 = _bsel_T[23]; // @[UserYanker.scala 92:55]
  wire  bsel_24 = _bsel_T[24]; // @[UserYanker.scala 92:55]
  wire  bsel_25 = _bsel_T[25]; // @[UserYanker.scala 92:55]
  wire  bsel_26 = _bsel_T[26]; // @[UserYanker.scala 92:55]
  wire  bsel_27 = _bsel_T[27]; // @[UserYanker.scala 92:55]
  wire  bsel_28 = _bsel_T[28]; // @[UserYanker.scala 92:55]
  wire  bsel_29 = _bsel_T[29]; // @[UserYanker.scala 92:55]
  wire  bsel_30 = _bsel_T[30]; // @[UserYanker.scala 92:55]
  wire  bsel_31 = _bsel_T[31]; // @[UserYanker.scala 92:55]
  wire  bsel_32 = _bsel_T[32]; // @[UserYanker.scala 92:55]
  wire  bsel_33 = _bsel_T[33]; // @[UserYanker.scala 92:55]
  wire  bsel_34 = _bsel_T[34]; // @[UserYanker.scala 92:55]
  wire  bsel_35 = _bsel_T[35]; // @[UserYanker.scala 92:55]
  wire  bsel_36 = _bsel_T[36]; // @[UserYanker.scala 92:55]
  wire  bsel_37 = _bsel_T[37]; // @[UserYanker.scala 92:55]
  wire  bsel_38 = _bsel_T[38]; // @[UserYanker.scala 92:55]
  wire  bsel_39 = _bsel_T[39]; // @[UserYanker.scala 92:55]
  wire  bsel_40 = _bsel_T[40]; // @[UserYanker.scala 92:55]
  wire  bsel_41 = _bsel_T[41]; // @[UserYanker.scala 92:55]
  wire  bsel_42 = _bsel_T[42]; // @[UserYanker.scala 92:55]
  wire  bsel_43 = _bsel_T[43]; // @[UserYanker.scala 92:55]
  wire  bsel_44 = _bsel_T[44]; // @[UserYanker.scala 92:55]
  wire  bsel_45 = _bsel_T[45]; // @[UserYanker.scala 92:55]
  wire  bsel_46 = _bsel_T[46]; // @[UserYanker.scala 92:55]
  wire  bsel_47 = _bsel_T[47]; // @[UserYanker.scala 92:55]
  wire  bsel_48 = _bsel_T[48]; // @[UserYanker.scala 92:55]
  wire  bsel_49 = _bsel_T[49]; // @[UserYanker.scala 92:55]
  wire  bsel_50 = _bsel_T[50]; // @[UserYanker.scala 92:55]
  wire  bsel_51 = _bsel_T[51]; // @[UserYanker.scala 92:55]
  wire  bsel_52 = _bsel_T[52]; // @[UserYanker.scala 92:55]
  wire  bsel_53 = _bsel_T[53]; // @[UserYanker.scala 92:55]
  wire  bsel_54 = _bsel_T[54]; // @[UserYanker.scala 92:55]
  wire  bsel_55 = _bsel_T[55]; // @[UserYanker.scala 92:55]
  wire  bsel_56 = _bsel_T[56]; // @[UserYanker.scala 92:55]
  wire  bsel_57 = _bsel_T[57]; // @[UserYanker.scala 92:55]
  wire  bsel_58 = _bsel_T[58]; // @[UserYanker.scala 92:55]
  wire  bsel_59 = _bsel_T[59]; // @[UserYanker.scala 92:55]
  wire  bsel_60 = _bsel_T[60]; // @[UserYanker.scala 92:55]
  wire  bsel_61 = _bsel_T[61]; // @[UserYanker.scala 92:55]
  wire  bsel_62 = _bsel_T[62]; // @[UserYanker.scala 92:55]
  wire  bsel_63 = _bsel_T[63]; // @[UserYanker.scala 92:55]
  Queue_33 Queue ( // @[UserYanker.scala 50:17]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_io_enq_bits_extra_id),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_io_deq_bits_extra_id)
  );
  Queue_33 Queue_1 ( // @[UserYanker.scala 50:17]
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_1_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_1_io_enq_bits_extra_id),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_1_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_1_io_deq_bits_extra_id)
  );
  Queue_35 Queue_2 ( // @[UserYanker.scala 50:17]
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_2_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_2_io_enq_bits_extra_id),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_2_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_2_io_deq_bits_extra_id)
  );
  Queue_35 Queue_3 ( // @[UserYanker.scala 50:17]
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_3_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_3_io_enq_bits_extra_id),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_3_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_3_io_deq_bits_extra_id)
  );
  Queue_35 Queue_4 ( // @[UserYanker.scala 50:17]
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_4_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_4_io_enq_bits_extra_id),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_4_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_4_io_deq_bits_extra_id)
  );
  Queue_35 Queue_5 ( // @[UserYanker.scala 50:17]
    .clock(Queue_5_clock),
    .reset(Queue_5_reset),
    .io_enq_ready(Queue_5_io_enq_ready),
    .io_enq_valid(Queue_5_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_5_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_5_io_enq_bits_extra_id),
    .io_deq_ready(Queue_5_io_deq_ready),
    .io_deq_valid(Queue_5_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_5_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_5_io_deq_bits_extra_id)
  );
  Queue_35 Queue_6 ( // @[UserYanker.scala 50:17]
    .clock(Queue_6_clock),
    .reset(Queue_6_reset),
    .io_enq_ready(Queue_6_io_enq_ready),
    .io_enq_valid(Queue_6_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_6_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_6_io_enq_bits_extra_id),
    .io_deq_ready(Queue_6_io_deq_ready),
    .io_deq_valid(Queue_6_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_6_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_6_io_deq_bits_extra_id)
  );
  Queue_35 Queue_7 ( // @[UserYanker.scala 50:17]
    .clock(Queue_7_clock),
    .reset(Queue_7_reset),
    .io_enq_ready(Queue_7_io_enq_ready),
    .io_enq_valid(Queue_7_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_7_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_7_io_enq_bits_extra_id),
    .io_deq_ready(Queue_7_io_deq_ready),
    .io_deq_valid(Queue_7_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_7_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_7_io_deq_bits_extra_id)
  );
  Queue_35 Queue_8 ( // @[UserYanker.scala 50:17]
    .clock(Queue_8_clock),
    .reset(Queue_8_reset),
    .io_enq_ready(Queue_8_io_enq_ready),
    .io_enq_valid(Queue_8_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_8_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_8_io_enq_bits_extra_id),
    .io_deq_ready(Queue_8_io_deq_ready),
    .io_deq_valid(Queue_8_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_8_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_8_io_deq_bits_extra_id)
  );
  Queue_35 Queue_9 ( // @[UserYanker.scala 50:17]
    .clock(Queue_9_clock),
    .reset(Queue_9_reset),
    .io_enq_ready(Queue_9_io_enq_ready),
    .io_enq_valid(Queue_9_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_9_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_9_io_enq_bits_extra_id),
    .io_deq_ready(Queue_9_io_deq_ready),
    .io_deq_valid(Queue_9_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_9_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_9_io_deq_bits_extra_id)
  );
  Queue_35 Queue_10 ( // @[UserYanker.scala 50:17]
    .clock(Queue_10_clock),
    .reset(Queue_10_reset),
    .io_enq_ready(Queue_10_io_enq_ready),
    .io_enq_valid(Queue_10_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_10_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_10_io_enq_bits_extra_id),
    .io_deq_ready(Queue_10_io_deq_ready),
    .io_deq_valid(Queue_10_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_10_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_10_io_deq_bits_extra_id)
  );
  Queue_35 Queue_11 ( // @[UserYanker.scala 50:17]
    .clock(Queue_11_clock),
    .reset(Queue_11_reset),
    .io_enq_ready(Queue_11_io_enq_ready),
    .io_enq_valid(Queue_11_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_11_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_11_io_enq_bits_extra_id),
    .io_deq_ready(Queue_11_io_deq_ready),
    .io_deq_valid(Queue_11_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_11_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_11_io_deq_bits_extra_id)
  );
  Queue_35 Queue_12 ( // @[UserYanker.scala 50:17]
    .clock(Queue_12_clock),
    .reset(Queue_12_reset),
    .io_enq_ready(Queue_12_io_enq_ready),
    .io_enq_valid(Queue_12_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_12_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_12_io_enq_bits_extra_id),
    .io_deq_ready(Queue_12_io_deq_ready),
    .io_deq_valid(Queue_12_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_12_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_12_io_deq_bits_extra_id)
  );
  Queue_35 Queue_13 ( // @[UserYanker.scala 50:17]
    .clock(Queue_13_clock),
    .reset(Queue_13_reset),
    .io_enq_ready(Queue_13_io_enq_ready),
    .io_enq_valid(Queue_13_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_13_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_13_io_enq_bits_extra_id),
    .io_deq_ready(Queue_13_io_deq_ready),
    .io_deq_valid(Queue_13_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_13_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_13_io_deq_bits_extra_id)
  );
  Queue_35 Queue_14 ( // @[UserYanker.scala 50:17]
    .clock(Queue_14_clock),
    .reset(Queue_14_reset),
    .io_enq_ready(Queue_14_io_enq_ready),
    .io_enq_valid(Queue_14_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_14_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_14_io_enq_bits_extra_id),
    .io_deq_ready(Queue_14_io_deq_ready),
    .io_deq_valid(Queue_14_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_14_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_14_io_deq_bits_extra_id)
  );
  Queue_35 Queue_15 ( // @[UserYanker.scala 50:17]
    .clock(Queue_15_clock),
    .reset(Queue_15_reset),
    .io_enq_ready(Queue_15_io_enq_ready),
    .io_enq_valid(Queue_15_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_15_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_15_io_enq_bits_extra_id),
    .io_deq_ready(Queue_15_io_deq_ready),
    .io_deq_valid(Queue_15_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_15_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_15_io_deq_bits_extra_id)
  );
  Queue_35 Queue_16 ( // @[UserYanker.scala 50:17]
    .clock(Queue_16_clock),
    .reset(Queue_16_reset),
    .io_enq_ready(Queue_16_io_enq_ready),
    .io_enq_valid(Queue_16_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_16_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_16_io_enq_bits_extra_id),
    .io_deq_ready(Queue_16_io_deq_ready),
    .io_deq_valid(Queue_16_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_16_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_16_io_deq_bits_extra_id)
  );
  Queue_35 Queue_17 ( // @[UserYanker.scala 50:17]
    .clock(Queue_17_clock),
    .reset(Queue_17_reset),
    .io_enq_ready(Queue_17_io_enq_ready),
    .io_enq_valid(Queue_17_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_17_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_17_io_enq_bits_extra_id),
    .io_deq_ready(Queue_17_io_deq_ready),
    .io_deq_valid(Queue_17_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_17_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_17_io_deq_bits_extra_id)
  );
  Queue_35 Queue_18 ( // @[UserYanker.scala 50:17]
    .clock(Queue_18_clock),
    .reset(Queue_18_reset),
    .io_enq_ready(Queue_18_io_enq_ready),
    .io_enq_valid(Queue_18_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_18_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_18_io_enq_bits_extra_id),
    .io_deq_ready(Queue_18_io_deq_ready),
    .io_deq_valid(Queue_18_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_18_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_18_io_deq_bits_extra_id)
  );
  Queue_35 Queue_19 ( // @[UserYanker.scala 50:17]
    .clock(Queue_19_clock),
    .reset(Queue_19_reset),
    .io_enq_ready(Queue_19_io_enq_ready),
    .io_enq_valid(Queue_19_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_19_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_19_io_enq_bits_extra_id),
    .io_deq_ready(Queue_19_io_deq_ready),
    .io_deq_valid(Queue_19_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_19_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_19_io_deq_bits_extra_id)
  );
  Queue_35 Queue_20 ( // @[UserYanker.scala 50:17]
    .clock(Queue_20_clock),
    .reset(Queue_20_reset),
    .io_enq_ready(Queue_20_io_enq_ready),
    .io_enq_valid(Queue_20_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_20_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_20_io_enq_bits_extra_id),
    .io_deq_ready(Queue_20_io_deq_ready),
    .io_deq_valid(Queue_20_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_20_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_20_io_deq_bits_extra_id)
  );
  Queue_35 Queue_21 ( // @[UserYanker.scala 50:17]
    .clock(Queue_21_clock),
    .reset(Queue_21_reset),
    .io_enq_ready(Queue_21_io_enq_ready),
    .io_enq_valid(Queue_21_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_21_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_21_io_enq_bits_extra_id),
    .io_deq_ready(Queue_21_io_deq_ready),
    .io_deq_valid(Queue_21_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_21_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_21_io_deq_bits_extra_id)
  );
  Queue_35 Queue_22 ( // @[UserYanker.scala 50:17]
    .clock(Queue_22_clock),
    .reset(Queue_22_reset),
    .io_enq_ready(Queue_22_io_enq_ready),
    .io_enq_valid(Queue_22_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_22_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_22_io_enq_bits_extra_id),
    .io_deq_ready(Queue_22_io_deq_ready),
    .io_deq_valid(Queue_22_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_22_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_22_io_deq_bits_extra_id)
  );
  Queue_35 Queue_23 ( // @[UserYanker.scala 50:17]
    .clock(Queue_23_clock),
    .reset(Queue_23_reset),
    .io_enq_ready(Queue_23_io_enq_ready),
    .io_enq_valid(Queue_23_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_23_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_23_io_enq_bits_extra_id),
    .io_deq_ready(Queue_23_io_deq_ready),
    .io_deq_valid(Queue_23_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_23_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_23_io_deq_bits_extra_id)
  );
  Queue_35 Queue_24 ( // @[UserYanker.scala 50:17]
    .clock(Queue_24_clock),
    .reset(Queue_24_reset),
    .io_enq_ready(Queue_24_io_enq_ready),
    .io_enq_valid(Queue_24_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_24_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_24_io_enq_bits_extra_id),
    .io_deq_ready(Queue_24_io_deq_ready),
    .io_deq_valid(Queue_24_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_24_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_24_io_deq_bits_extra_id)
  );
  Queue_35 Queue_25 ( // @[UserYanker.scala 50:17]
    .clock(Queue_25_clock),
    .reset(Queue_25_reset),
    .io_enq_ready(Queue_25_io_enq_ready),
    .io_enq_valid(Queue_25_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_25_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_25_io_enq_bits_extra_id),
    .io_deq_ready(Queue_25_io_deq_ready),
    .io_deq_valid(Queue_25_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_25_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_25_io_deq_bits_extra_id)
  );
  Queue_35 Queue_26 ( // @[UserYanker.scala 50:17]
    .clock(Queue_26_clock),
    .reset(Queue_26_reset),
    .io_enq_ready(Queue_26_io_enq_ready),
    .io_enq_valid(Queue_26_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_26_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_26_io_enq_bits_extra_id),
    .io_deq_ready(Queue_26_io_deq_ready),
    .io_deq_valid(Queue_26_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_26_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_26_io_deq_bits_extra_id)
  );
  Queue_35 Queue_27 ( // @[UserYanker.scala 50:17]
    .clock(Queue_27_clock),
    .reset(Queue_27_reset),
    .io_enq_ready(Queue_27_io_enq_ready),
    .io_enq_valid(Queue_27_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_27_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_27_io_enq_bits_extra_id),
    .io_deq_ready(Queue_27_io_deq_ready),
    .io_deq_valid(Queue_27_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_27_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_27_io_deq_bits_extra_id)
  );
  Queue_35 Queue_28 ( // @[UserYanker.scala 50:17]
    .clock(Queue_28_clock),
    .reset(Queue_28_reset),
    .io_enq_ready(Queue_28_io_enq_ready),
    .io_enq_valid(Queue_28_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_28_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_28_io_enq_bits_extra_id),
    .io_deq_ready(Queue_28_io_deq_ready),
    .io_deq_valid(Queue_28_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_28_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_28_io_deq_bits_extra_id)
  );
  Queue_35 Queue_29 ( // @[UserYanker.scala 50:17]
    .clock(Queue_29_clock),
    .reset(Queue_29_reset),
    .io_enq_ready(Queue_29_io_enq_ready),
    .io_enq_valid(Queue_29_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_29_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_29_io_enq_bits_extra_id),
    .io_deq_ready(Queue_29_io_deq_ready),
    .io_deq_valid(Queue_29_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_29_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_29_io_deq_bits_extra_id)
  );
  Queue_35 Queue_30 ( // @[UserYanker.scala 50:17]
    .clock(Queue_30_clock),
    .reset(Queue_30_reset),
    .io_enq_ready(Queue_30_io_enq_ready),
    .io_enq_valid(Queue_30_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_30_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_30_io_enq_bits_extra_id),
    .io_deq_ready(Queue_30_io_deq_ready),
    .io_deq_valid(Queue_30_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_30_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_30_io_deq_bits_extra_id)
  );
  Queue_35 Queue_31 ( // @[UserYanker.scala 50:17]
    .clock(Queue_31_clock),
    .reset(Queue_31_reset),
    .io_enq_ready(Queue_31_io_enq_ready),
    .io_enq_valid(Queue_31_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_31_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_31_io_enq_bits_extra_id),
    .io_deq_ready(Queue_31_io_deq_ready),
    .io_deq_valid(Queue_31_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_31_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_31_io_deq_bits_extra_id)
  );
  Queue_35 Queue_32 ( // @[UserYanker.scala 50:17]
    .clock(Queue_32_clock),
    .reset(Queue_32_reset),
    .io_enq_ready(Queue_32_io_enq_ready),
    .io_enq_valid(Queue_32_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_32_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_32_io_enq_bits_extra_id),
    .io_deq_ready(Queue_32_io_deq_ready),
    .io_deq_valid(Queue_32_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_32_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_32_io_deq_bits_extra_id)
  );
  Queue_35 Queue_33 ( // @[UserYanker.scala 50:17]
    .clock(Queue_33_clock),
    .reset(Queue_33_reset),
    .io_enq_ready(Queue_33_io_enq_ready),
    .io_enq_valid(Queue_33_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_33_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_33_io_enq_bits_extra_id),
    .io_deq_ready(Queue_33_io_deq_ready),
    .io_deq_valid(Queue_33_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_33_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_33_io_deq_bits_extra_id)
  );
  Queue_35 Queue_34 ( // @[UserYanker.scala 50:17]
    .clock(Queue_34_clock),
    .reset(Queue_34_reset),
    .io_enq_ready(Queue_34_io_enq_ready),
    .io_enq_valid(Queue_34_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_34_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_34_io_enq_bits_extra_id),
    .io_deq_ready(Queue_34_io_deq_ready),
    .io_deq_valid(Queue_34_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_34_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_34_io_deq_bits_extra_id)
  );
  Queue_35 Queue_35 ( // @[UserYanker.scala 50:17]
    .clock(Queue_35_clock),
    .reset(Queue_35_reset),
    .io_enq_ready(Queue_35_io_enq_ready),
    .io_enq_valid(Queue_35_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_35_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_35_io_enq_bits_extra_id),
    .io_deq_ready(Queue_35_io_deq_ready),
    .io_deq_valid(Queue_35_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_35_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_35_io_deq_bits_extra_id)
  );
  Queue_35 Queue_36 ( // @[UserYanker.scala 50:17]
    .clock(Queue_36_clock),
    .reset(Queue_36_reset),
    .io_enq_ready(Queue_36_io_enq_ready),
    .io_enq_valid(Queue_36_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_36_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_36_io_enq_bits_extra_id),
    .io_deq_ready(Queue_36_io_deq_ready),
    .io_deq_valid(Queue_36_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_36_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_36_io_deq_bits_extra_id)
  );
  Queue_35 Queue_37 ( // @[UserYanker.scala 50:17]
    .clock(Queue_37_clock),
    .reset(Queue_37_reset),
    .io_enq_ready(Queue_37_io_enq_ready),
    .io_enq_valid(Queue_37_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_37_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_37_io_enq_bits_extra_id),
    .io_deq_ready(Queue_37_io_deq_ready),
    .io_deq_valid(Queue_37_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_37_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_37_io_deq_bits_extra_id)
  );
  Queue_35 Queue_38 ( // @[UserYanker.scala 50:17]
    .clock(Queue_38_clock),
    .reset(Queue_38_reset),
    .io_enq_ready(Queue_38_io_enq_ready),
    .io_enq_valid(Queue_38_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_38_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_38_io_enq_bits_extra_id),
    .io_deq_ready(Queue_38_io_deq_ready),
    .io_deq_valid(Queue_38_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_38_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_38_io_deq_bits_extra_id)
  );
  Queue_35 Queue_39 ( // @[UserYanker.scala 50:17]
    .clock(Queue_39_clock),
    .reset(Queue_39_reset),
    .io_enq_ready(Queue_39_io_enq_ready),
    .io_enq_valid(Queue_39_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_39_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_39_io_enq_bits_extra_id),
    .io_deq_ready(Queue_39_io_deq_ready),
    .io_deq_valid(Queue_39_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_39_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_39_io_deq_bits_extra_id)
  );
  Queue_35 Queue_40 ( // @[UserYanker.scala 50:17]
    .clock(Queue_40_clock),
    .reset(Queue_40_reset),
    .io_enq_ready(Queue_40_io_enq_ready),
    .io_enq_valid(Queue_40_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_40_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_40_io_enq_bits_extra_id),
    .io_deq_ready(Queue_40_io_deq_ready),
    .io_deq_valid(Queue_40_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_40_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_40_io_deq_bits_extra_id)
  );
  Queue_35 Queue_41 ( // @[UserYanker.scala 50:17]
    .clock(Queue_41_clock),
    .reset(Queue_41_reset),
    .io_enq_ready(Queue_41_io_enq_ready),
    .io_enq_valid(Queue_41_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_41_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_41_io_enq_bits_extra_id),
    .io_deq_ready(Queue_41_io_deq_ready),
    .io_deq_valid(Queue_41_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_41_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_41_io_deq_bits_extra_id)
  );
  Queue_35 Queue_42 ( // @[UserYanker.scala 50:17]
    .clock(Queue_42_clock),
    .reset(Queue_42_reset),
    .io_enq_ready(Queue_42_io_enq_ready),
    .io_enq_valid(Queue_42_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_42_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_42_io_enq_bits_extra_id),
    .io_deq_ready(Queue_42_io_deq_ready),
    .io_deq_valid(Queue_42_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_42_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_42_io_deq_bits_extra_id)
  );
  Queue_35 Queue_43 ( // @[UserYanker.scala 50:17]
    .clock(Queue_43_clock),
    .reset(Queue_43_reset),
    .io_enq_ready(Queue_43_io_enq_ready),
    .io_enq_valid(Queue_43_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_43_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_43_io_enq_bits_extra_id),
    .io_deq_ready(Queue_43_io_deq_ready),
    .io_deq_valid(Queue_43_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_43_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_43_io_deq_bits_extra_id)
  );
  Queue_35 Queue_44 ( // @[UserYanker.scala 50:17]
    .clock(Queue_44_clock),
    .reset(Queue_44_reset),
    .io_enq_ready(Queue_44_io_enq_ready),
    .io_enq_valid(Queue_44_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_44_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_44_io_enq_bits_extra_id),
    .io_deq_ready(Queue_44_io_deq_ready),
    .io_deq_valid(Queue_44_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_44_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_44_io_deq_bits_extra_id)
  );
  Queue_35 Queue_45 ( // @[UserYanker.scala 50:17]
    .clock(Queue_45_clock),
    .reset(Queue_45_reset),
    .io_enq_ready(Queue_45_io_enq_ready),
    .io_enq_valid(Queue_45_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_45_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_45_io_enq_bits_extra_id),
    .io_deq_ready(Queue_45_io_deq_ready),
    .io_deq_valid(Queue_45_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_45_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_45_io_deq_bits_extra_id)
  );
  Queue_35 Queue_46 ( // @[UserYanker.scala 50:17]
    .clock(Queue_46_clock),
    .reset(Queue_46_reset),
    .io_enq_ready(Queue_46_io_enq_ready),
    .io_enq_valid(Queue_46_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_46_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_46_io_enq_bits_extra_id),
    .io_deq_ready(Queue_46_io_deq_ready),
    .io_deq_valid(Queue_46_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_46_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_46_io_deq_bits_extra_id)
  );
  Queue_35 Queue_47 ( // @[UserYanker.scala 50:17]
    .clock(Queue_47_clock),
    .reset(Queue_47_reset),
    .io_enq_ready(Queue_47_io_enq_ready),
    .io_enq_valid(Queue_47_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_47_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_47_io_enq_bits_extra_id),
    .io_deq_ready(Queue_47_io_deq_ready),
    .io_deq_valid(Queue_47_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_47_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_47_io_deq_bits_extra_id)
  );
  Queue_35 Queue_48 ( // @[UserYanker.scala 50:17]
    .clock(Queue_48_clock),
    .reset(Queue_48_reset),
    .io_enq_ready(Queue_48_io_enq_ready),
    .io_enq_valid(Queue_48_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_48_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_48_io_enq_bits_extra_id),
    .io_deq_ready(Queue_48_io_deq_ready),
    .io_deq_valid(Queue_48_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_48_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_48_io_deq_bits_extra_id)
  );
  Queue_35 Queue_49 ( // @[UserYanker.scala 50:17]
    .clock(Queue_49_clock),
    .reset(Queue_49_reset),
    .io_enq_ready(Queue_49_io_enq_ready),
    .io_enq_valid(Queue_49_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_49_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_49_io_enq_bits_extra_id),
    .io_deq_ready(Queue_49_io_deq_ready),
    .io_deq_valid(Queue_49_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_49_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_49_io_deq_bits_extra_id)
  );
  Queue_35 Queue_50 ( // @[UserYanker.scala 50:17]
    .clock(Queue_50_clock),
    .reset(Queue_50_reset),
    .io_enq_ready(Queue_50_io_enq_ready),
    .io_enq_valid(Queue_50_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_50_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_50_io_enq_bits_extra_id),
    .io_deq_ready(Queue_50_io_deq_ready),
    .io_deq_valid(Queue_50_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_50_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_50_io_deq_bits_extra_id)
  );
  Queue_35 Queue_51 ( // @[UserYanker.scala 50:17]
    .clock(Queue_51_clock),
    .reset(Queue_51_reset),
    .io_enq_ready(Queue_51_io_enq_ready),
    .io_enq_valid(Queue_51_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_51_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_51_io_enq_bits_extra_id),
    .io_deq_ready(Queue_51_io_deq_ready),
    .io_deq_valid(Queue_51_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_51_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_51_io_deq_bits_extra_id)
  );
  Queue_35 Queue_52 ( // @[UserYanker.scala 50:17]
    .clock(Queue_52_clock),
    .reset(Queue_52_reset),
    .io_enq_ready(Queue_52_io_enq_ready),
    .io_enq_valid(Queue_52_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_52_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_52_io_enq_bits_extra_id),
    .io_deq_ready(Queue_52_io_deq_ready),
    .io_deq_valid(Queue_52_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_52_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_52_io_deq_bits_extra_id)
  );
  Queue_35 Queue_53 ( // @[UserYanker.scala 50:17]
    .clock(Queue_53_clock),
    .reset(Queue_53_reset),
    .io_enq_ready(Queue_53_io_enq_ready),
    .io_enq_valid(Queue_53_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_53_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_53_io_enq_bits_extra_id),
    .io_deq_ready(Queue_53_io_deq_ready),
    .io_deq_valid(Queue_53_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_53_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_53_io_deq_bits_extra_id)
  );
  Queue_35 Queue_54 ( // @[UserYanker.scala 50:17]
    .clock(Queue_54_clock),
    .reset(Queue_54_reset),
    .io_enq_ready(Queue_54_io_enq_ready),
    .io_enq_valid(Queue_54_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_54_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_54_io_enq_bits_extra_id),
    .io_deq_ready(Queue_54_io_deq_ready),
    .io_deq_valid(Queue_54_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_54_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_54_io_deq_bits_extra_id)
  );
  Queue_35 Queue_55 ( // @[UserYanker.scala 50:17]
    .clock(Queue_55_clock),
    .reset(Queue_55_reset),
    .io_enq_ready(Queue_55_io_enq_ready),
    .io_enq_valid(Queue_55_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_55_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_55_io_enq_bits_extra_id),
    .io_deq_ready(Queue_55_io_deq_ready),
    .io_deq_valid(Queue_55_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_55_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_55_io_deq_bits_extra_id)
  );
  Queue_35 Queue_56 ( // @[UserYanker.scala 50:17]
    .clock(Queue_56_clock),
    .reset(Queue_56_reset),
    .io_enq_ready(Queue_56_io_enq_ready),
    .io_enq_valid(Queue_56_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_56_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_56_io_enq_bits_extra_id),
    .io_deq_ready(Queue_56_io_deq_ready),
    .io_deq_valid(Queue_56_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_56_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_56_io_deq_bits_extra_id)
  );
  Queue_35 Queue_57 ( // @[UserYanker.scala 50:17]
    .clock(Queue_57_clock),
    .reset(Queue_57_reset),
    .io_enq_ready(Queue_57_io_enq_ready),
    .io_enq_valid(Queue_57_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_57_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_57_io_enq_bits_extra_id),
    .io_deq_ready(Queue_57_io_deq_ready),
    .io_deq_valid(Queue_57_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_57_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_57_io_deq_bits_extra_id)
  );
  Queue_35 Queue_58 ( // @[UserYanker.scala 50:17]
    .clock(Queue_58_clock),
    .reset(Queue_58_reset),
    .io_enq_ready(Queue_58_io_enq_ready),
    .io_enq_valid(Queue_58_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_58_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_58_io_enq_bits_extra_id),
    .io_deq_ready(Queue_58_io_deq_ready),
    .io_deq_valid(Queue_58_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_58_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_58_io_deq_bits_extra_id)
  );
  Queue_35 Queue_59 ( // @[UserYanker.scala 50:17]
    .clock(Queue_59_clock),
    .reset(Queue_59_reset),
    .io_enq_ready(Queue_59_io_enq_ready),
    .io_enq_valid(Queue_59_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_59_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_59_io_enq_bits_extra_id),
    .io_deq_ready(Queue_59_io_deq_ready),
    .io_deq_valid(Queue_59_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_59_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_59_io_deq_bits_extra_id)
  );
  Queue_35 Queue_60 ( // @[UserYanker.scala 50:17]
    .clock(Queue_60_clock),
    .reset(Queue_60_reset),
    .io_enq_ready(Queue_60_io_enq_ready),
    .io_enq_valid(Queue_60_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_60_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_60_io_enq_bits_extra_id),
    .io_deq_ready(Queue_60_io_deq_ready),
    .io_deq_valid(Queue_60_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_60_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_60_io_deq_bits_extra_id)
  );
  Queue_35 Queue_61 ( // @[UserYanker.scala 50:17]
    .clock(Queue_61_clock),
    .reset(Queue_61_reset),
    .io_enq_ready(Queue_61_io_enq_ready),
    .io_enq_valid(Queue_61_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_61_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_61_io_enq_bits_extra_id),
    .io_deq_ready(Queue_61_io_deq_ready),
    .io_deq_valid(Queue_61_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_61_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_61_io_deq_bits_extra_id)
  );
  Queue_35 Queue_62 ( // @[UserYanker.scala 50:17]
    .clock(Queue_62_clock),
    .reset(Queue_62_reset),
    .io_enq_ready(Queue_62_io_enq_ready),
    .io_enq_valid(Queue_62_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_62_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_62_io_enq_bits_extra_id),
    .io_deq_ready(Queue_62_io_deq_ready),
    .io_deq_valid(Queue_62_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_62_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_62_io_deq_bits_extra_id)
  );
  Queue_35 Queue_63 ( // @[UserYanker.scala 50:17]
    .clock(Queue_63_clock),
    .reset(Queue_63_reset),
    .io_enq_ready(Queue_63_io_enq_ready),
    .io_enq_valid(Queue_63_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_63_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_63_io_enq_bits_extra_id),
    .io_deq_ready(Queue_63_io_deq_ready),
    .io_deq_valid(Queue_63_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_63_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_63_io_deq_bits_extra_id)
  );
  Queue_33 Queue_64 ( // @[UserYanker.scala 50:17]
    .clock(Queue_64_clock),
    .reset(Queue_64_reset),
    .io_enq_ready(Queue_64_io_enq_ready),
    .io_enq_valid(Queue_64_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_64_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_64_io_enq_bits_extra_id),
    .io_deq_ready(Queue_64_io_deq_ready),
    .io_deq_valid(Queue_64_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_64_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_64_io_deq_bits_extra_id)
  );
  Queue_33 Queue_65 ( // @[UserYanker.scala 50:17]
    .clock(Queue_65_clock),
    .reset(Queue_65_reset),
    .io_enq_ready(Queue_65_io_enq_ready),
    .io_enq_valid(Queue_65_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_65_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_65_io_enq_bits_extra_id),
    .io_deq_ready(Queue_65_io_deq_ready),
    .io_deq_valid(Queue_65_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_65_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_65_io_deq_bits_extra_id)
  );
  Queue_35 Queue_66 ( // @[UserYanker.scala 50:17]
    .clock(Queue_66_clock),
    .reset(Queue_66_reset),
    .io_enq_ready(Queue_66_io_enq_ready),
    .io_enq_valid(Queue_66_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_66_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_66_io_enq_bits_extra_id),
    .io_deq_ready(Queue_66_io_deq_ready),
    .io_deq_valid(Queue_66_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_66_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_66_io_deq_bits_extra_id)
  );
  Queue_35 Queue_67 ( // @[UserYanker.scala 50:17]
    .clock(Queue_67_clock),
    .reset(Queue_67_reset),
    .io_enq_ready(Queue_67_io_enq_ready),
    .io_enq_valid(Queue_67_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_67_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_67_io_enq_bits_extra_id),
    .io_deq_ready(Queue_67_io_deq_ready),
    .io_deq_valid(Queue_67_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_67_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_67_io_deq_bits_extra_id)
  );
  Queue_35 Queue_68 ( // @[UserYanker.scala 50:17]
    .clock(Queue_68_clock),
    .reset(Queue_68_reset),
    .io_enq_ready(Queue_68_io_enq_ready),
    .io_enq_valid(Queue_68_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_68_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_68_io_enq_bits_extra_id),
    .io_deq_ready(Queue_68_io_deq_ready),
    .io_deq_valid(Queue_68_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_68_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_68_io_deq_bits_extra_id)
  );
  Queue_35 Queue_69 ( // @[UserYanker.scala 50:17]
    .clock(Queue_69_clock),
    .reset(Queue_69_reset),
    .io_enq_ready(Queue_69_io_enq_ready),
    .io_enq_valid(Queue_69_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_69_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_69_io_enq_bits_extra_id),
    .io_deq_ready(Queue_69_io_deq_ready),
    .io_deq_valid(Queue_69_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_69_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_69_io_deq_bits_extra_id)
  );
  Queue_35 Queue_70 ( // @[UserYanker.scala 50:17]
    .clock(Queue_70_clock),
    .reset(Queue_70_reset),
    .io_enq_ready(Queue_70_io_enq_ready),
    .io_enq_valid(Queue_70_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_70_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_70_io_enq_bits_extra_id),
    .io_deq_ready(Queue_70_io_deq_ready),
    .io_deq_valid(Queue_70_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_70_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_70_io_deq_bits_extra_id)
  );
  Queue_35 Queue_71 ( // @[UserYanker.scala 50:17]
    .clock(Queue_71_clock),
    .reset(Queue_71_reset),
    .io_enq_ready(Queue_71_io_enq_ready),
    .io_enq_valid(Queue_71_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_71_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_71_io_enq_bits_extra_id),
    .io_deq_ready(Queue_71_io_deq_ready),
    .io_deq_valid(Queue_71_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_71_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_71_io_deq_bits_extra_id)
  );
  Queue_35 Queue_72 ( // @[UserYanker.scala 50:17]
    .clock(Queue_72_clock),
    .reset(Queue_72_reset),
    .io_enq_ready(Queue_72_io_enq_ready),
    .io_enq_valid(Queue_72_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_72_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_72_io_enq_bits_extra_id),
    .io_deq_ready(Queue_72_io_deq_ready),
    .io_deq_valid(Queue_72_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_72_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_72_io_deq_bits_extra_id)
  );
  Queue_35 Queue_73 ( // @[UserYanker.scala 50:17]
    .clock(Queue_73_clock),
    .reset(Queue_73_reset),
    .io_enq_ready(Queue_73_io_enq_ready),
    .io_enq_valid(Queue_73_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_73_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_73_io_enq_bits_extra_id),
    .io_deq_ready(Queue_73_io_deq_ready),
    .io_deq_valid(Queue_73_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_73_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_73_io_deq_bits_extra_id)
  );
  Queue_35 Queue_74 ( // @[UserYanker.scala 50:17]
    .clock(Queue_74_clock),
    .reset(Queue_74_reset),
    .io_enq_ready(Queue_74_io_enq_ready),
    .io_enq_valid(Queue_74_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_74_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_74_io_enq_bits_extra_id),
    .io_deq_ready(Queue_74_io_deq_ready),
    .io_deq_valid(Queue_74_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_74_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_74_io_deq_bits_extra_id)
  );
  Queue_35 Queue_75 ( // @[UserYanker.scala 50:17]
    .clock(Queue_75_clock),
    .reset(Queue_75_reset),
    .io_enq_ready(Queue_75_io_enq_ready),
    .io_enq_valid(Queue_75_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_75_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_75_io_enq_bits_extra_id),
    .io_deq_ready(Queue_75_io_deq_ready),
    .io_deq_valid(Queue_75_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_75_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_75_io_deq_bits_extra_id)
  );
  Queue_35 Queue_76 ( // @[UserYanker.scala 50:17]
    .clock(Queue_76_clock),
    .reset(Queue_76_reset),
    .io_enq_ready(Queue_76_io_enq_ready),
    .io_enq_valid(Queue_76_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_76_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_76_io_enq_bits_extra_id),
    .io_deq_ready(Queue_76_io_deq_ready),
    .io_deq_valid(Queue_76_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_76_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_76_io_deq_bits_extra_id)
  );
  Queue_35 Queue_77 ( // @[UserYanker.scala 50:17]
    .clock(Queue_77_clock),
    .reset(Queue_77_reset),
    .io_enq_ready(Queue_77_io_enq_ready),
    .io_enq_valid(Queue_77_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_77_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_77_io_enq_bits_extra_id),
    .io_deq_ready(Queue_77_io_deq_ready),
    .io_deq_valid(Queue_77_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_77_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_77_io_deq_bits_extra_id)
  );
  Queue_35 Queue_78 ( // @[UserYanker.scala 50:17]
    .clock(Queue_78_clock),
    .reset(Queue_78_reset),
    .io_enq_ready(Queue_78_io_enq_ready),
    .io_enq_valid(Queue_78_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_78_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_78_io_enq_bits_extra_id),
    .io_deq_ready(Queue_78_io_deq_ready),
    .io_deq_valid(Queue_78_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_78_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_78_io_deq_bits_extra_id)
  );
  Queue_35 Queue_79 ( // @[UserYanker.scala 50:17]
    .clock(Queue_79_clock),
    .reset(Queue_79_reset),
    .io_enq_ready(Queue_79_io_enq_ready),
    .io_enq_valid(Queue_79_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_79_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_79_io_enq_bits_extra_id),
    .io_deq_ready(Queue_79_io_deq_ready),
    .io_deq_valid(Queue_79_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_79_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_79_io_deq_bits_extra_id)
  );
  Queue_35 Queue_80 ( // @[UserYanker.scala 50:17]
    .clock(Queue_80_clock),
    .reset(Queue_80_reset),
    .io_enq_ready(Queue_80_io_enq_ready),
    .io_enq_valid(Queue_80_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_80_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_80_io_enq_bits_extra_id),
    .io_deq_ready(Queue_80_io_deq_ready),
    .io_deq_valid(Queue_80_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_80_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_80_io_deq_bits_extra_id)
  );
  Queue_35 Queue_81 ( // @[UserYanker.scala 50:17]
    .clock(Queue_81_clock),
    .reset(Queue_81_reset),
    .io_enq_ready(Queue_81_io_enq_ready),
    .io_enq_valid(Queue_81_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_81_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_81_io_enq_bits_extra_id),
    .io_deq_ready(Queue_81_io_deq_ready),
    .io_deq_valid(Queue_81_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_81_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_81_io_deq_bits_extra_id)
  );
  Queue_35 Queue_82 ( // @[UserYanker.scala 50:17]
    .clock(Queue_82_clock),
    .reset(Queue_82_reset),
    .io_enq_ready(Queue_82_io_enq_ready),
    .io_enq_valid(Queue_82_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_82_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_82_io_enq_bits_extra_id),
    .io_deq_ready(Queue_82_io_deq_ready),
    .io_deq_valid(Queue_82_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_82_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_82_io_deq_bits_extra_id)
  );
  Queue_35 Queue_83 ( // @[UserYanker.scala 50:17]
    .clock(Queue_83_clock),
    .reset(Queue_83_reset),
    .io_enq_ready(Queue_83_io_enq_ready),
    .io_enq_valid(Queue_83_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_83_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_83_io_enq_bits_extra_id),
    .io_deq_ready(Queue_83_io_deq_ready),
    .io_deq_valid(Queue_83_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_83_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_83_io_deq_bits_extra_id)
  );
  Queue_35 Queue_84 ( // @[UserYanker.scala 50:17]
    .clock(Queue_84_clock),
    .reset(Queue_84_reset),
    .io_enq_ready(Queue_84_io_enq_ready),
    .io_enq_valid(Queue_84_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_84_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_84_io_enq_bits_extra_id),
    .io_deq_ready(Queue_84_io_deq_ready),
    .io_deq_valid(Queue_84_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_84_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_84_io_deq_bits_extra_id)
  );
  Queue_35 Queue_85 ( // @[UserYanker.scala 50:17]
    .clock(Queue_85_clock),
    .reset(Queue_85_reset),
    .io_enq_ready(Queue_85_io_enq_ready),
    .io_enq_valid(Queue_85_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_85_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_85_io_enq_bits_extra_id),
    .io_deq_ready(Queue_85_io_deq_ready),
    .io_deq_valid(Queue_85_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_85_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_85_io_deq_bits_extra_id)
  );
  Queue_35 Queue_86 ( // @[UserYanker.scala 50:17]
    .clock(Queue_86_clock),
    .reset(Queue_86_reset),
    .io_enq_ready(Queue_86_io_enq_ready),
    .io_enq_valid(Queue_86_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_86_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_86_io_enq_bits_extra_id),
    .io_deq_ready(Queue_86_io_deq_ready),
    .io_deq_valid(Queue_86_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_86_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_86_io_deq_bits_extra_id)
  );
  Queue_35 Queue_87 ( // @[UserYanker.scala 50:17]
    .clock(Queue_87_clock),
    .reset(Queue_87_reset),
    .io_enq_ready(Queue_87_io_enq_ready),
    .io_enq_valid(Queue_87_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_87_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_87_io_enq_bits_extra_id),
    .io_deq_ready(Queue_87_io_deq_ready),
    .io_deq_valid(Queue_87_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_87_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_87_io_deq_bits_extra_id)
  );
  Queue_35 Queue_88 ( // @[UserYanker.scala 50:17]
    .clock(Queue_88_clock),
    .reset(Queue_88_reset),
    .io_enq_ready(Queue_88_io_enq_ready),
    .io_enq_valid(Queue_88_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_88_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_88_io_enq_bits_extra_id),
    .io_deq_ready(Queue_88_io_deq_ready),
    .io_deq_valid(Queue_88_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_88_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_88_io_deq_bits_extra_id)
  );
  Queue_35 Queue_89 ( // @[UserYanker.scala 50:17]
    .clock(Queue_89_clock),
    .reset(Queue_89_reset),
    .io_enq_ready(Queue_89_io_enq_ready),
    .io_enq_valid(Queue_89_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_89_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_89_io_enq_bits_extra_id),
    .io_deq_ready(Queue_89_io_deq_ready),
    .io_deq_valid(Queue_89_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_89_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_89_io_deq_bits_extra_id)
  );
  Queue_35 Queue_90 ( // @[UserYanker.scala 50:17]
    .clock(Queue_90_clock),
    .reset(Queue_90_reset),
    .io_enq_ready(Queue_90_io_enq_ready),
    .io_enq_valid(Queue_90_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_90_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_90_io_enq_bits_extra_id),
    .io_deq_ready(Queue_90_io_deq_ready),
    .io_deq_valid(Queue_90_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_90_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_90_io_deq_bits_extra_id)
  );
  Queue_35 Queue_91 ( // @[UserYanker.scala 50:17]
    .clock(Queue_91_clock),
    .reset(Queue_91_reset),
    .io_enq_ready(Queue_91_io_enq_ready),
    .io_enq_valid(Queue_91_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_91_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_91_io_enq_bits_extra_id),
    .io_deq_ready(Queue_91_io_deq_ready),
    .io_deq_valid(Queue_91_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_91_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_91_io_deq_bits_extra_id)
  );
  Queue_35 Queue_92 ( // @[UserYanker.scala 50:17]
    .clock(Queue_92_clock),
    .reset(Queue_92_reset),
    .io_enq_ready(Queue_92_io_enq_ready),
    .io_enq_valid(Queue_92_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_92_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_92_io_enq_bits_extra_id),
    .io_deq_ready(Queue_92_io_deq_ready),
    .io_deq_valid(Queue_92_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_92_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_92_io_deq_bits_extra_id)
  );
  Queue_35 Queue_93 ( // @[UserYanker.scala 50:17]
    .clock(Queue_93_clock),
    .reset(Queue_93_reset),
    .io_enq_ready(Queue_93_io_enq_ready),
    .io_enq_valid(Queue_93_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_93_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_93_io_enq_bits_extra_id),
    .io_deq_ready(Queue_93_io_deq_ready),
    .io_deq_valid(Queue_93_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_93_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_93_io_deq_bits_extra_id)
  );
  Queue_35 Queue_94 ( // @[UserYanker.scala 50:17]
    .clock(Queue_94_clock),
    .reset(Queue_94_reset),
    .io_enq_ready(Queue_94_io_enq_ready),
    .io_enq_valid(Queue_94_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_94_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_94_io_enq_bits_extra_id),
    .io_deq_ready(Queue_94_io_deq_ready),
    .io_deq_valid(Queue_94_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_94_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_94_io_deq_bits_extra_id)
  );
  Queue_35 Queue_95 ( // @[UserYanker.scala 50:17]
    .clock(Queue_95_clock),
    .reset(Queue_95_reset),
    .io_enq_ready(Queue_95_io_enq_ready),
    .io_enq_valid(Queue_95_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_95_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_95_io_enq_bits_extra_id),
    .io_deq_ready(Queue_95_io_deq_ready),
    .io_deq_valid(Queue_95_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_95_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_95_io_deq_bits_extra_id)
  );
  Queue_35 Queue_96 ( // @[UserYanker.scala 50:17]
    .clock(Queue_96_clock),
    .reset(Queue_96_reset),
    .io_enq_ready(Queue_96_io_enq_ready),
    .io_enq_valid(Queue_96_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_96_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_96_io_enq_bits_extra_id),
    .io_deq_ready(Queue_96_io_deq_ready),
    .io_deq_valid(Queue_96_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_96_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_96_io_deq_bits_extra_id)
  );
  Queue_35 Queue_97 ( // @[UserYanker.scala 50:17]
    .clock(Queue_97_clock),
    .reset(Queue_97_reset),
    .io_enq_ready(Queue_97_io_enq_ready),
    .io_enq_valid(Queue_97_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_97_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_97_io_enq_bits_extra_id),
    .io_deq_ready(Queue_97_io_deq_ready),
    .io_deq_valid(Queue_97_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_97_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_97_io_deq_bits_extra_id)
  );
  Queue_35 Queue_98 ( // @[UserYanker.scala 50:17]
    .clock(Queue_98_clock),
    .reset(Queue_98_reset),
    .io_enq_ready(Queue_98_io_enq_ready),
    .io_enq_valid(Queue_98_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_98_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_98_io_enq_bits_extra_id),
    .io_deq_ready(Queue_98_io_deq_ready),
    .io_deq_valid(Queue_98_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_98_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_98_io_deq_bits_extra_id)
  );
  Queue_35 Queue_99 ( // @[UserYanker.scala 50:17]
    .clock(Queue_99_clock),
    .reset(Queue_99_reset),
    .io_enq_ready(Queue_99_io_enq_ready),
    .io_enq_valid(Queue_99_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_99_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_99_io_enq_bits_extra_id),
    .io_deq_ready(Queue_99_io_deq_ready),
    .io_deq_valid(Queue_99_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_99_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_99_io_deq_bits_extra_id)
  );
  Queue_35 Queue_100 ( // @[UserYanker.scala 50:17]
    .clock(Queue_100_clock),
    .reset(Queue_100_reset),
    .io_enq_ready(Queue_100_io_enq_ready),
    .io_enq_valid(Queue_100_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_100_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_100_io_enq_bits_extra_id),
    .io_deq_ready(Queue_100_io_deq_ready),
    .io_deq_valid(Queue_100_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_100_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_100_io_deq_bits_extra_id)
  );
  Queue_35 Queue_101 ( // @[UserYanker.scala 50:17]
    .clock(Queue_101_clock),
    .reset(Queue_101_reset),
    .io_enq_ready(Queue_101_io_enq_ready),
    .io_enq_valid(Queue_101_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_101_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_101_io_enq_bits_extra_id),
    .io_deq_ready(Queue_101_io_deq_ready),
    .io_deq_valid(Queue_101_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_101_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_101_io_deq_bits_extra_id)
  );
  Queue_35 Queue_102 ( // @[UserYanker.scala 50:17]
    .clock(Queue_102_clock),
    .reset(Queue_102_reset),
    .io_enq_ready(Queue_102_io_enq_ready),
    .io_enq_valid(Queue_102_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_102_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_102_io_enq_bits_extra_id),
    .io_deq_ready(Queue_102_io_deq_ready),
    .io_deq_valid(Queue_102_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_102_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_102_io_deq_bits_extra_id)
  );
  Queue_35 Queue_103 ( // @[UserYanker.scala 50:17]
    .clock(Queue_103_clock),
    .reset(Queue_103_reset),
    .io_enq_ready(Queue_103_io_enq_ready),
    .io_enq_valid(Queue_103_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_103_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_103_io_enq_bits_extra_id),
    .io_deq_ready(Queue_103_io_deq_ready),
    .io_deq_valid(Queue_103_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_103_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_103_io_deq_bits_extra_id)
  );
  Queue_35 Queue_104 ( // @[UserYanker.scala 50:17]
    .clock(Queue_104_clock),
    .reset(Queue_104_reset),
    .io_enq_ready(Queue_104_io_enq_ready),
    .io_enq_valid(Queue_104_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_104_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_104_io_enq_bits_extra_id),
    .io_deq_ready(Queue_104_io_deq_ready),
    .io_deq_valid(Queue_104_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_104_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_104_io_deq_bits_extra_id)
  );
  Queue_35 Queue_105 ( // @[UserYanker.scala 50:17]
    .clock(Queue_105_clock),
    .reset(Queue_105_reset),
    .io_enq_ready(Queue_105_io_enq_ready),
    .io_enq_valid(Queue_105_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_105_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_105_io_enq_bits_extra_id),
    .io_deq_ready(Queue_105_io_deq_ready),
    .io_deq_valid(Queue_105_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_105_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_105_io_deq_bits_extra_id)
  );
  Queue_35 Queue_106 ( // @[UserYanker.scala 50:17]
    .clock(Queue_106_clock),
    .reset(Queue_106_reset),
    .io_enq_ready(Queue_106_io_enq_ready),
    .io_enq_valid(Queue_106_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_106_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_106_io_enq_bits_extra_id),
    .io_deq_ready(Queue_106_io_deq_ready),
    .io_deq_valid(Queue_106_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_106_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_106_io_deq_bits_extra_id)
  );
  Queue_35 Queue_107 ( // @[UserYanker.scala 50:17]
    .clock(Queue_107_clock),
    .reset(Queue_107_reset),
    .io_enq_ready(Queue_107_io_enq_ready),
    .io_enq_valid(Queue_107_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_107_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_107_io_enq_bits_extra_id),
    .io_deq_ready(Queue_107_io_deq_ready),
    .io_deq_valid(Queue_107_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_107_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_107_io_deq_bits_extra_id)
  );
  Queue_35 Queue_108 ( // @[UserYanker.scala 50:17]
    .clock(Queue_108_clock),
    .reset(Queue_108_reset),
    .io_enq_ready(Queue_108_io_enq_ready),
    .io_enq_valid(Queue_108_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_108_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_108_io_enq_bits_extra_id),
    .io_deq_ready(Queue_108_io_deq_ready),
    .io_deq_valid(Queue_108_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_108_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_108_io_deq_bits_extra_id)
  );
  Queue_35 Queue_109 ( // @[UserYanker.scala 50:17]
    .clock(Queue_109_clock),
    .reset(Queue_109_reset),
    .io_enq_ready(Queue_109_io_enq_ready),
    .io_enq_valid(Queue_109_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_109_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_109_io_enq_bits_extra_id),
    .io_deq_ready(Queue_109_io_deq_ready),
    .io_deq_valid(Queue_109_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_109_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_109_io_deq_bits_extra_id)
  );
  Queue_35 Queue_110 ( // @[UserYanker.scala 50:17]
    .clock(Queue_110_clock),
    .reset(Queue_110_reset),
    .io_enq_ready(Queue_110_io_enq_ready),
    .io_enq_valid(Queue_110_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_110_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_110_io_enq_bits_extra_id),
    .io_deq_ready(Queue_110_io_deq_ready),
    .io_deq_valid(Queue_110_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_110_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_110_io_deq_bits_extra_id)
  );
  Queue_35 Queue_111 ( // @[UserYanker.scala 50:17]
    .clock(Queue_111_clock),
    .reset(Queue_111_reset),
    .io_enq_ready(Queue_111_io_enq_ready),
    .io_enq_valid(Queue_111_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_111_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_111_io_enq_bits_extra_id),
    .io_deq_ready(Queue_111_io_deq_ready),
    .io_deq_valid(Queue_111_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_111_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_111_io_deq_bits_extra_id)
  );
  Queue_35 Queue_112 ( // @[UserYanker.scala 50:17]
    .clock(Queue_112_clock),
    .reset(Queue_112_reset),
    .io_enq_ready(Queue_112_io_enq_ready),
    .io_enq_valid(Queue_112_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_112_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_112_io_enq_bits_extra_id),
    .io_deq_ready(Queue_112_io_deq_ready),
    .io_deq_valid(Queue_112_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_112_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_112_io_deq_bits_extra_id)
  );
  Queue_35 Queue_113 ( // @[UserYanker.scala 50:17]
    .clock(Queue_113_clock),
    .reset(Queue_113_reset),
    .io_enq_ready(Queue_113_io_enq_ready),
    .io_enq_valid(Queue_113_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_113_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_113_io_enq_bits_extra_id),
    .io_deq_ready(Queue_113_io_deq_ready),
    .io_deq_valid(Queue_113_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_113_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_113_io_deq_bits_extra_id)
  );
  Queue_35 Queue_114 ( // @[UserYanker.scala 50:17]
    .clock(Queue_114_clock),
    .reset(Queue_114_reset),
    .io_enq_ready(Queue_114_io_enq_ready),
    .io_enq_valid(Queue_114_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_114_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_114_io_enq_bits_extra_id),
    .io_deq_ready(Queue_114_io_deq_ready),
    .io_deq_valid(Queue_114_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_114_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_114_io_deq_bits_extra_id)
  );
  Queue_35 Queue_115 ( // @[UserYanker.scala 50:17]
    .clock(Queue_115_clock),
    .reset(Queue_115_reset),
    .io_enq_ready(Queue_115_io_enq_ready),
    .io_enq_valid(Queue_115_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_115_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_115_io_enq_bits_extra_id),
    .io_deq_ready(Queue_115_io_deq_ready),
    .io_deq_valid(Queue_115_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_115_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_115_io_deq_bits_extra_id)
  );
  Queue_35 Queue_116 ( // @[UserYanker.scala 50:17]
    .clock(Queue_116_clock),
    .reset(Queue_116_reset),
    .io_enq_ready(Queue_116_io_enq_ready),
    .io_enq_valid(Queue_116_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_116_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_116_io_enq_bits_extra_id),
    .io_deq_ready(Queue_116_io_deq_ready),
    .io_deq_valid(Queue_116_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_116_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_116_io_deq_bits_extra_id)
  );
  Queue_35 Queue_117 ( // @[UserYanker.scala 50:17]
    .clock(Queue_117_clock),
    .reset(Queue_117_reset),
    .io_enq_ready(Queue_117_io_enq_ready),
    .io_enq_valid(Queue_117_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_117_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_117_io_enq_bits_extra_id),
    .io_deq_ready(Queue_117_io_deq_ready),
    .io_deq_valid(Queue_117_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_117_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_117_io_deq_bits_extra_id)
  );
  Queue_35 Queue_118 ( // @[UserYanker.scala 50:17]
    .clock(Queue_118_clock),
    .reset(Queue_118_reset),
    .io_enq_ready(Queue_118_io_enq_ready),
    .io_enq_valid(Queue_118_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_118_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_118_io_enq_bits_extra_id),
    .io_deq_ready(Queue_118_io_deq_ready),
    .io_deq_valid(Queue_118_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_118_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_118_io_deq_bits_extra_id)
  );
  Queue_35 Queue_119 ( // @[UserYanker.scala 50:17]
    .clock(Queue_119_clock),
    .reset(Queue_119_reset),
    .io_enq_ready(Queue_119_io_enq_ready),
    .io_enq_valid(Queue_119_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_119_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_119_io_enq_bits_extra_id),
    .io_deq_ready(Queue_119_io_deq_ready),
    .io_deq_valid(Queue_119_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_119_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_119_io_deq_bits_extra_id)
  );
  Queue_35 Queue_120 ( // @[UserYanker.scala 50:17]
    .clock(Queue_120_clock),
    .reset(Queue_120_reset),
    .io_enq_ready(Queue_120_io_enq_ready),
    .io_enq_valid(Queue_120_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_120_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_120_io_enq_bits_extra_id),
    .io_deq_ready(Queue_120_io_deq_ready),
    .io_deq_valid(Queue_120_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_120_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_120_io_deq_bits_extra_id)
  );
  Queue_35 Queue_121 ( // @[UserYanker.scala 50:17]
    .clock(Queue_121_clock),
    .reset(Queue_121_reset),
    .io_enq_ready(Queue_121_io_enq_ready),
    .io_enq_valid(Queue_121_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_121_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_121_io_enq_bits_extra_id),
    .io_deq_ready(Queue_121_io_deq_ready),
    .io_deq_valid(Queue_121_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_121_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_121_io_deq_bits_extra_id)
  );
  Queue_35 Queue_122 ( // @[UserYanker.scala 50:17]
    .clock(Queue_122_clock),
    .reset(Queue_122_reset),
    .io_enq_ready(Queue_122_io_enq_ready),
    .io_enq_valid(Queue_122_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_122_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_122_io_enq_bits_extra_id),
    .io_deq_ready(Queue_122_io_deq_ready),
    .io_deq_valid(Queue_122_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_122_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_122_io_deq_bits_extra_id)
  );
  Queue_35 Queue_123 ( // @[UserYanker.scala 50:17]
    .clock(Queue_123_clock),
    .reset(Queue_123_reset),
    .io_enq_ready(Queue_123_io_enq_ready),
    .io_enq_valid(Queue_123_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_123_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_123_io_enq_bits_extra_id),
    .io_deq_ready(Queue_123_io_deq_ready),
    .io_deq_valid(Queue_123_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_123_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_123_io_deq_bits_extra_id)
  );
  Queue_35 Queue_124 ( // @[UserYanker.scala 50:17]
    .clock(Queue_124_clock),
    .reset(Queue_124_reset),
    .io_enq_ready(Queue_124_io_enq_ready),
    .io_enq_valid(Queue_124_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_124_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_124_io_enq_bits_extra_id),
    .io_deq_ready(Queue_124_io_deq_ready),
    .io_deq_valid(Queue_124_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_124_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_124_io_deq_bits_extra_id)
  );
  Queue_35 Queue_125 ( // @[UserYanker.scala 50:17]
    .clock(Queue_125_clock),
    .reset(Queue_125_reset),
    .io_enq_ready(Queue_125_io_enq_ready),
    .io_enq_valid(Queue_125_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_125_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_125_io_enq_bits_extra_id),
    .io_deq_ready(Queue_125_io_deq_ready),
    .io_deq_valid(Queue_125_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_125_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_125_io_deq_bits_extra_id)
  );
  Queue_35 Queue_126 ( // @[UserYanker.scala 50:17]
    .clock(Queue_126_clock),
    .reset(Queue_126_reset),
    .io_enq_ready(Queue_126_io_enq_ready),
    .io_enq_valid(Queue_126_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_126_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_126_io_enq_bits_extra_id),
    .io_deq_ready(Queue_126_io_deq_ready),
    .io_deq_valid(Queue_126_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_126_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_126_io_deq_bits_extra_id)
  );
  Queue_35 Queue_127 ( // @[UserYanker.scala 50:17]
    .clock(Queue_127_clock),
    .reset(Queue_127_reset),
    .io_enq_ready(Queue_127_io_enq_ready),
    .io_enq_valid(Queue_127_io_enq_valid),
    .io_enq_bits_tl_state_source(Queue_127_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(Queue_127_io_enq_bits_extra_id),
    .io_deq_ready(Queue_127_io_deq_ready),
    .io_deq_valid(Queue_127_io_deq_valid),
    .io_deq_bits_tl_state_source(Queue_127_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(Queue_127_io_deq_bits_extra_id)
  );
  assign auto_in_aw_ready = auto_out_aw_ready & _GEN_383; // @[UserYanker.scala 80:36]
  assign auto_in_w_ready = auto_out_w_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_b_valid = auto_out_b_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_b_bits_id = auto_out_b_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_b_bits_echo_tl_state_source = 6'h3f == auto_out_b_bits_id ? _b_bits_WIRE_63_tl_state_source : _GEN_574; // @[BundleMap.scala 247:{19,19}]
  assign auto_in_b_bits_echo_extra_id = 6'h3f == auto_out_b_bits_id ? _b_bits_WIRE_63_extra_id : _GEN_510; // @[BundleMap.scala 247:{19,19}]
  assign auto_in_ar_ready = auto_out_ar_ready & _GEN_63; // @[UserYanker.scala 59:36]
  assign auto_in_r_valid = auto_out_r_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_bits_id = auto_out_r_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_bits_echo_tl_state_source = 6'h3f == auto_out_r_bits_id ? _r_bits_WIRE_63_tl_state_source : _GEN_254; // @[BundleMap.scala 247:{19,19}]
  assign auto_in_r_bits_echo_extra_id = 6'h3f == auto_out_r_bits_id ? _r_bits_WIRE_63_extra_id : _GEN_190; // @[BundleMap.scala 247:{19,19}]
  assign auto_in_r_bits_last = auto_out_r_bits_last; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_out_aw_valid = auto_in_aw_valid & _GEN_383; // @[UserYanker.scala 81:36]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_len = auto_in_aw_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_size = auto_in_aw_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_burst = auto_in_aw_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_lock = auto_in_aw_bits_lock; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_cache = auto_in_aw_bits_cache; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_prot = auto_in_aw_bits_prot; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_qos = auto_in_aw_bits_qos; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_w_valid = auto_in_w_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_w_bits_strb = auto_in_w_bits_strb; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_b_ready = auto_in_b_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_valid = auto_in_ar_valid & _GEN_63; // @[UserYanker.scala 60:36]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_len = auto_in_ar_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_burst = auto_in_ar_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_lock = auto_in_ar_bits_lock; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_cache = auto_in_ar_bits_cache; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_prot = auto_in_ar_bits_prot; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_qos = auto_in_ar_bits_qos; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_r_ready = auto_in_r_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_0; // @[UserYanker.scala 74:53]
  assign Queue_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_0 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_1; // @[UserYanker.scala 74:53]
  assign Queue_1_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_1_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_1_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_1 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign Queue_2_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_2; // @[UserYanker.scala 74:53]
  assign Queue_2_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_2_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_2_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_2 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign Queue_3_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_3; // @[UserYanker.scala 74:53]
  assign Queue_3_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_3_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_3_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_3 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_4_clock = clock;
  assign Queue_4_reset = reset;
  assign Queue_4_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_4; // @[UserYanker.scala 74:53]
  assign Queue_4_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_4_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_4_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_4 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_5_clock = clock;
  assign Queue_5_reset = reset;
  assign Queue_5_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_5; // @[UserYanker.scala 74:53]
  assign Queue_5_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_5_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_5_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_5 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_6_clock = clock;
  assign Queue_6_reset = reset;
  assign Queue_6_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_6; // @[UserYanker.scala 74:53]
  assign Queue_6_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_6_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_6_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_6 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_7_clock = clock;
  assign Queue_7_reset = reset;
  assign Queue_7_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_7; // @[UserYanker.scala 74:53]
  assign Queue_7_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_7_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_7_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_7 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_8_clock = clock;
  assign Queue_8_reset = reset;
  assign Queue_8_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_8; // @[UserYanker.scala 74:53]
  assign Queue_8_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_8_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_8_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_8 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_9_clock = clock;
  assign Queue_9_reset = reset;
  assign Queue_9_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_9; // @[UserYanker.scala 74:53]
  assign Queue_9_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_9_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_9_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_9 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_10_clock = clock;
  assign Queue_10_reset = reset;
  assign Queue_10_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_10; // @[UserYanker.scala 74:53]
  assign Queue_10_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_10_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_10_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_10 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_11_clock = clock;
  assign Queue_11_reset = reset;
  assign Queue_11_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_11; // @[UserYanker.scala 74:53]
  assign Queue_11_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_11_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_11_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_11 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_12_clock = clock;
  assign Queue_12_reset = reset;
  assign Queue_12_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_12; // @[UserYanker.scala 74:53]
  assign Queue_12_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_12_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_12_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_12 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_13_clock = clock;
  assign Queue_13_reset = reset;
  assign Queue_13_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_13; // @[UserYanker.scala 74:53]
  assign Queue_13_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_13_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_13_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_13 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_14_clock = clock;
  assign Queue_14_reset = reset;
  assign Queue_14_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_14; // @[UserYanker.scala 74:53]
  assign Queue_14_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_14_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_14_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_14 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_15_clock = clock;
  assign Queue_15_reset = reset;
  assign Queue_15_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_15; // @[UserYanker.scala 74:53]
  assign Queue_15_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_15_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_15_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_15 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_16_clock = clock;
  assign Queue_16_reset = reset;
  assign Queue_16_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_16; // @[UserYanker.scala 74:53]
  assign Queue_16_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_16_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_16_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_16 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_17_clock = clock;
  assign Queue_17_reset = reset;
  assign Queue_17_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_17; // @[UserYanker.scala 74:53]
  assign Queue_17_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_17_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_17_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_17 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_18_clock = clock;
  assign Queue_18_reset = reset;
  assign Queue_18_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_18; // @[UserYanker.scala 74:53]
  assign Queue_18_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_18_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_18_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_18 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_19_clock = clock;
  assign Queue_19_reset = reset;
  assign Queue_19_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_19; // @[UserYanker.scala 74:53]
  assign Queue_19_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_19_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_19_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_19 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_20_clock = clock;
  assign Queue_20_reset = reset;
  assign Queue_20_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_20; // @[UserYanker.scala 74:53]
  assign Queue_20_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_20_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_20_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_20 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_21_clock = clock;
  assign Queue_21_reset = reset;
  assign Queue_21_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_21; // @[UserYanker.scala 74:53]
  assign Queue_21_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_21_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_21_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_21 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_22_clock = clock;
  assign Queue_22_reset = reset;
  assign Queue_22_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_22; // @[UserYanker.scala 74:53]
  assign Queue_22_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_22_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_22_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_22 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_23_clock = clock;
  assign Queue_23_reset = reset;
  assign Queue_23_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_23; // @[UserYanker.scala 74:53]
  assign Queue_23_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_23_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_23_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_23 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_24_clock = clock;
  assign Queue_24_reset = reset;
  assign Queue_24_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_24; // @[UserYanker.scala 74:53]
  assign Queue_24_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_24_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_24_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_24 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_25_clock = clock;
  assign Queue_25_reset = reset;
  assign Queue_25_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_25; // @[UserYanker.scala 74:53]
  assign Queue_25_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_25_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_25_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_25 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_26_clock = clock;
  assign Queue_26_reset = reset;
  assign Queue_26_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_26; // @[UserYanker.scala 74:53]
  assign Queue_26_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_26_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_26_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_26 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_27_clock = clock;
  assign Queue_27_reset = reset;
  assign Queue_27_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_27; // @[UserYanker.scala 74:53]
  assign Queue_27_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_27_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_27_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_27 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_28_clock = clock;
  assign Queue_28_reset = reset;
  assign Queue_28_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_28; // @[UserYanker.scala 74:53]
  assign Queue_28_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_28_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_28_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_28 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_29_clock = clock;
  assign Queue_29_reset = reset;
  assign Queue_29_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_29; // @[UserYanker.scala 74:53]
  assign Queue_29_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_29_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_29_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_29 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_30_clock = clock;
  assign Queue_30_reset = reset;
  assign Queue_30_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_30; // @[UserYanker.scala 74:53]
  assign Queue_30_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_30_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_30_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_30 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_31_clock = clock;
  assign Queue_31_reset = reset;
  assign Queue_31_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_31; // @[UserYanker.scala 74:53]
  assign Queue_31_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_31_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_31_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_31 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_32_clock = clock;
  assign Queue_32_reset = reset;
  assign Queue_32_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_32; // @[UserYanker.scala 74:53]
  assign Queue_32_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_32_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_32_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_32 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_33_clock = clock;
  assign Queue_33_reset = reset;
  assign Queue_33_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_33; // @[UserYanker.scala 74:53]
  assign Queue_33_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_33_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_33_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_33 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_34_clock = clock;
  assign Queue_34_reset = reset;
  assign Queue_34_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_34; // @[UserYanker.scala 74:53]
  assign Queue_34_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_34_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_34_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_34 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_35_clock = clock;
  assign Queue_35_reset = reset;
  assign Queue_35_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_35; // @[UserYanker.scala 74:53]
  assign Queue_35_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_35_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_35_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_35 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_36_clock = clock;
  assign Queue_36_reset = reset;
  assign Queue_36_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_36; // @[UserYanker.scala 74:53]
  assign Queue_36_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_36_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_36_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_36 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_37_clock = clock;
  assign Queue_37_reset = reset;
  assign Queue_37_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_37; // @[UserYanker.scala 74:53]
  assign Queue_37_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_37_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_37_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_37 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_38_clock = clock;
  assign Queue_38_reset = reset;
  assign Queue_38_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_38; // @[UserYanker.scala 74:53]
  assign Queue_38_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_38_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_38_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_38 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_39_clock = clock;
  assign Queue_39_reset = reset;
  assign Queue_39_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_39; // @[UserYanker.scala 74:53]
  assign Queue_39_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_39_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_39_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_39 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_40_clock = clock;
  assign Queue_40_reset = reset;
  assign Queue_40_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_40; // @[UserYanker.scala 74:53]
  assign Queue_40_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_40_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_40_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_40 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_41_clock = clock;
  assign Queue_41_reset = reset;
  assign Queue_41_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_41; // @[UserYanker.scala 74:53]
  assign Queue_41_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_41_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_41_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_41 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_42_clock = clock;
  assign Queue_42_reset = reset;
  assign Queue_42_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_42; // @[UserYanker.scala 74:53]
  assign Queue_42_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_42_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_42_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_42 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_43_clock = clock;
  assign Queue_43_reset = reset;
  assign Queue_43_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_43; // @[UserYanker.scala 74:53]
  assign Queue_43_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_43_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_43_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_43 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_44_clock = clock;
  assign Queue_44_reset = reset;
  assign Queue_44_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_44; // @[UserYanker.scala 74:53]
  assign Queue_44_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_44_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_44_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_44 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_45_clock = clock;
  assign Queue_45_reset = reset;
  assign Queue_45_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_45; // @[UserYanker.scala 74:53]
  assign Queue_45_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_45_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_45_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_45 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_46_clock = clock;
  assign Queue_46_reset = reset;
  assign Queue_46_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_46; // @[UserYanker.scala 74:53]
  assign Queue_46_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_46_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_46_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_46 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_47_clock = clock;
  assign Queue_47_reset = reset;
  assign Queue_47_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_47; // @[UserYanker.scala 74:53]
  assign Queue_47_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_47_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_47_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_47 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_48_clock = clock;
  assign Queue_48_reset = reset;
  assign Queue_48_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_48; // @[UserYanker.scala 74:53]
  assign Queue_48_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_48_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_48_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_48 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_49_clock = clock;
  assign Queue_49_reset = reset;
  assign Queue_49_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_49; // @[UserYanker.scala 74:53]
  assign Queue_49_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_49_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_49_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_49 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_50_clock = clock;
  assign Queue_50_reset = reset;
  assign Queue_50_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_50; // @[UserYanker.scala 74:53]
  assign Queue_50_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_50_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_50_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_50 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_51_clock = clock;
  assign Queue_51_reset = reset;
  assign Queue_51_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_51; // @[UserYanker.scala 74:53]
  assign Queue_51_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_51_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_51_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_51 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_52_clock = clock;
  assign Queue_52_reset = reset;
  assign Queue_52_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_52; // @[UserYanker.scala 74:53]
  assign Queue_52_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_52_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_52_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_52 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_53_clock = clock;
  assign Queue_53_reset = reset;
  assign Queue_53_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_53; // @[UserYanker.scala 74:53]
  assign Queue_53_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_53_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_53_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_53 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_54_clock = clock;
  assign Queue_54_reset = reset;
  assign Queue_54_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_54; // @[UserYanker.scala 74:53]
  assign Queue_54_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_54_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_54_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_54 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_55_clock = clock;
  assign Queue_55_reset = reset;
  assign Queue_55_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_55; // @[UserYanker.scala 74:53]
  assign Queue_55_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_55_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_55_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_55 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_56_clock = clock;
  assign Queue_56_reset = reset;
  assign Queue_56_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_56; // @[UserYanker.scala 74:53]
  assign Queue_56_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_56_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_56_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_56 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_57_clock = clock;
  assign Queue_57_reset = reset;
  assign Queue_57_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_57; // @[UserYanker.scala 74:53]
  assign Queue_57_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_57_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_57_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_57 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_58_clock = clock;
  assign Queue_58_reset = reset;
  assign Queue_58_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_58; // @[UserYanker.scala 74:53]
  assign Queue_58_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_58_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_58_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_58 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_59_clock = clock;
  assign Queue_59_reset = reset;
  assign Queue_59_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_59; // @[UserYanker.scala 74:53]
  assign Queue_59_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_59_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_59_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_59 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_60_clock = clock;
  assign Queue_60_reset = reset;
  assign Queue_60_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_60; // @[UserYanker.scala 74:53]
  assign Queue_60_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_60_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_60_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_60 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_61_clock = clock;
  assign Queue_61_reset = reset;
  assign Queue_61_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_61; // @[UserYanker.scala 74:53]
  assign Queue_61_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_61_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_61_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_61 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_62_clock = clock;
  assign Queue_62_reset = reset;
  assign Queue_62_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_62; // @[UserYanker.scala 74:53]
  assign Queue_62_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_62_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_62_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_62 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_63_clock = clock;
  assign Queue_63_reset = reset;
  assign Queue_63_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_63; // @[UserYanker.scala 74:53]
  assign Queue_63_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_63_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_63_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_63 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_64_clock = clock;
  assign Queue_64_reset = reset;
  assign Queue_64_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_0; // @[UserYanker.scala 95:53]
  assign Queue_64_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_64_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_64_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_0; // @[UserYanker.scala 94:53]
  assign Queue_65_clock = clock;
  assign Queue_65_reset = reset;
  assign Queue_65_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_1; // @[UserYanker.scala 95:53]
  assign Queue_65_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_65_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_65_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_1; // @[UserYanker.scala 94:53]
  assign Queue_66_clock = clock;
  assign Queue_66_reset = reset;
  assign Queue_66_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_2; // @[UserYanker.scala 95:53]
  assign Queue_66_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_66_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_66_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_2; // @[UserYanker.scala 94:53]
  assign Queue_67_clock = clock;
  assign Queue_67_reset = reset;
  assign Queue_67_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_3; // @[UserYanker.scala 95:53]
  assign Queue_67_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_67_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_67_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_3; // @[UserYanker.scala 94:53]
  assign Queue_68_clock = clock;
  assign Queue_68_reset = reset;
  assign Queue_68_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_4; // @[UserYanker.scala 95:53]
  assign Queue_68_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_68_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_68_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_4; // @[UserYanker.scala 94:53]
  assign Queue_69_clock = clock;
  assign Queue_69_reset = reset;
  assign Queue_69_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_5; // @[UserYanker.scala 95:53]
  assign Queue_69_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_69_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_69_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_5; // @[UserYanker.scala 94:53]
  assign Queue_70_clock = clock;
  assign Queue_70_reset = reset;
  assign Queue_70_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_6; // @[UserYanker.scala 95:53]
  assign Queue_70_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_70_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_70_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_6; // @[UserYanker.scala 94:53]
  assign Queue_71_clock = clock;
  assign Queue_71_reset = reset;
  assign Queue_71_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_7; // @[UserYanker.scala 95:53]
  assign Queue_71_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_71_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_71_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_7; // @[UserYanker.scala 94:53]
  assign Queue_72_clock = clock;
  assign Queue_72_reset = reset;
  assign Queue_72_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_8; // @[UserYanker.scala 95:53]
  assign Queue_72_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_72_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_72_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_8; // @[UserYanker.scala 94:53]
  assign Queue_73_clock = clock;
  assign Queue_73_reset = reset;
  assign Queue_73_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_9; // @[UserYanker.scala 95:53]
  assign Queue_73_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_73_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_73_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_9; // @[UserYanker.scala 94:53]
  assign Queue_74_clock = clock;
  assign Queue_74_reset = reset;
  assign Queue_74_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_10; // @[UserYanker.scala 95:53]
  assign Queue_74_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_74_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_74_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_10; // @[UserYanker.scala 94:53]
  assign Queue_75_clock = clock;
  assign Queue_75_reset = reset;
  assign Queue_75_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_11; // @[UserYanker.scala 95:53]
  assign Queue_75_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_75_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_75_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_11; // @[UserYanker.scala 94:53]
  assign Queue_76_clock = clock;
  assign Queue_76_reset = reset;
  assign Queue_76_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_12; // @[UserYanker.scala 95:53]
  assign Queue_76_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_76_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_76_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_12; // @[UserYanker.scala 94:53]
  assign Queue_77_clock = clock;
  assign Queue_77_reset = reset;
  assign Queue_77_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_13; // @[UserYanker.scala 95:53]
  assign Queue_77_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_77_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_77_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_13; // @[UserYanker.scala 94:53]
  assign Queue_78_clock = clock;
  assign Queue_78_reset = reset;
  assign Queue_78_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_14; // @[UserYanker.scala 95:53]
  assign Queue_78_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_78_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_78_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_14; // @[UserYanker.scala 94:53]
  assign Queue_79_clock = clock;
  assign Queue_79_reset = reset;
  assign Queue_79_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_15; // @[UserYanker.scala 95:53]
  assign Queue_79_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_79_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_79_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_15; // @[UserYanker.scala 94:53]
  assign Queue_80_clock = clock;
  assign Queue_80_reset = reset;
  assign Queue_80_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_16; // @[UserYanker.scala 95:53]
  assign Queue_80_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_80_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_80_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_16; // @[UserYanker.scala 94:53]
  assign Queue_81_clock = clock;
  assign Queue_81_reset = reset;
  assign Queue_81_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_17; // @[UserYanker.scala 95:53]
  assign Queue_81_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_81_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_81_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_17; // @[UserYanker.scala 94:53]
  assign Queue_82_clock = clock;
  assign Queue_82_reset = reset;
  assign Queue_82_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_18; // @[UserYanker.scala 95:53]
  assign Queue_82_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_82_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_82_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_18; // @[UserYanker.scala 94:53]
  assign Queue_83_clock = clock;
  assign Queue_83_reset = reset;
  assign Queue_83_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_19; // @[UserYanker.scala 95:53]
  assign Queue_83_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_83_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_83_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_19; // @[UserYanker.scala 94:53]
  assign Queue_84_clock = clock;
  assign Queue_84_reset = reset;
  assign Queue_84_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_20; // @[UserYanker.scala 95:53]
  assign Queue_84_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_84_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_84_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_20; // @[UserYanker.scala 94:53]
  assign Queue_85_clock = clock;
  assign Queue_85_reset = reset;
  assign Queue_85_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_21; // @[UserYanker.scala 95:53]
  assign Queue_85_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_85_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_85_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_21; // @[UserYanker.scala 94:53]
  assign Queue_86_clock = clock;
  assign Queue_86_reset = reset;
  assign Queue_86_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_22; // @[UserYanker.scala 95:53]
  assign Queue_86_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_86_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_86_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_22; // @[UserYanker.scala 94:53]
  assign Queue_87_clock = clock;
  assign Queue_87_reset = reset;
  assign Queue_87_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_23; // @[UserYanker.scala 95:53]
  assign Queue_87_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_87_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_87_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_23; // @[UserYanker.scala 94:53]
  assign Queue_88_clock = clock;
  assign Queue_88_reset = reset;
  assign Queue_88_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_24; // @[UserYanker.scala 95:53]
  assign Queue_88_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_88_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_88_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_24; // @[UserYanker.scala 94:53]
  assign Queue_89_clock = clock;
  assign Queue_89_reset = reset;
  assign Queue_89_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_25; // @[UserYanker.scala 95:53]
  assign Queue_89_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_89_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_89_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_25; // @[UserYanker.scala 94:53]
  assign Queue_90_clock = clock;
  assign Queue_90_reset = reset;
  assign Queue_90_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_26; // @[UserYanker.scala 95:53]
  assign Queue_90_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_90_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_90_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_26; // @[UserYanker.scala 94:53]
  assign Queue_91_clock = clock;
  assign Queue_91_reset = reset;
  assign Queue_91_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_27; // @[UserYanker.scala 95:53]
  assign Queue_91_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_91_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_91_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_27; // @[UserYanker.scala 94:53]
  assign Queue_92_clock = clock;
  assign Queue_92_reset = reset;
  assign Queue_92_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_28; // @[UserYanker.scala 95:53]
  assign Queue_92_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_92_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_92_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_28; // @[UserYanker.scala 94:53]
  assign Queue_93_clock = clock;
  assign Queue_93_reset = reset;
  assign Queue_93_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_29; // @[UserYanker.scala 95:53]
  assign Queue_93_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_93_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_93_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_29; // @[UserYanker.scala 94:53]
  assign Queue_94_clock = clock;
  assign Queue_94_reset = reset;
  assign Queue_94_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_30; // @[UserYanker.scala 95:53]
  assign Queue_94_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_94_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_94_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_30; // @[UserYanker.scala 94:53]
  assign Queue_95_clock = clock;
  assign Queue_95_reset = reset;
  assign Queue_95_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_31; // @[UserYanker.scala 95:53]
  assign Queue_95_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_95_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_95_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_31; // @[UserYanker.scala 94:53]
  assign Queue_96_clock = clock;
  assign Queue_96_reset = reset;
  assign Queue_96_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_32; // @[UserYanker.scala 95:53]
  assign Queue_96_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_96_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_96_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_32; // @[UserYanker.scala 94:53]
  assign Queue_97_clock = clock;
  assign Queue_97_reset = reset;
  assign Queue_97_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_33; // @[UserYanker.scala 95:53]
  assign Queue_97_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_97_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_97_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_33; // @[UserYanker.scala 94:53]
  assign Queue_98_clock = clock;
  assign Queue_98_reset = reset;
  assign Queue_98_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_34; // @[UserYanker.scala 95:53]
  assign Queue_98_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_98_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_98_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_34; // @[UserYanker.scala 94:53]
  assign Queue_99_clock = clock;
  assign Queue_99_reset = reset;
  assign Queue_99_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_35; // @[UserYanker.scala 95:53]
  assign Queue_99_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_99_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_99_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_35; // @[UserYanker.scala 94:53]
  assign Queue_100_clock = clock;
  assign Queue_100_reset = reset;
  assign Queue_100_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_36; // @[UserYanker.scala 95:53]
  assign Queue_100_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_100_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_100_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_36; // @[UserYanker.scala 94:53]
  assign Queue_101_clock = clock;
  assign Queue_101_reset = reset;
  assign Queue_101_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_37; // @[UserYanker.scala 95:53]
  assign Queue_101_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_101_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_101_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_37; // @[UserYanker.scala 94:53]
  assign Queue_102_clock = clock;
  assign Queue_102_reset = reset;
  assign Queue_102_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_38; // @[UserYanker.scala 95:53]
  assign Queue_102_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_102_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_102_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_38; // @[UserYanker.scala 94:53]
  assign Queue_103_clock = clock;
  assign Queue_103_reset = reset;
  assign Queue_103_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_39; // @[UserYanker.scala 95:53]
  assign Queue_103_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_103_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_103_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_39; // @[UserYanker.scala 94:53]
  assign Queue_104_clock = clock;
  assign Queue_104_reset = reset;
  assign Queue_104_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_40; // @[UserYanker.scala 95:53]
  assign Queue_104_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_104_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_104_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_40; // @[UserYanker.scala 94:53]
  assign Queue_105_clock = clock;
  assign Queue_105_reset = reset;
  assign Queue_105_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_41; // @[UserYanker.scala 95:53]
  assign Queue_105_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_105_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_105_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_41; // @[UserYanker.scala 94:53]
  assign Queue_106_clock = clock;
  assign Queue_106_reset = reset;
  assign Queue_106_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_42; // @[UserYanker.scala 95:53]
  assign Queue_106_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_106_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_106_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_42; // @[UserYanker.scala 94:53]
  assign Queue_107_clock = clock;
  assign Queue_107_reset = reset;
  assign Queue_107_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_43; // @[UserYanker.scala 95:53]
  assign Queue_107_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_107_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_107_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_43; // @[UserYanker.scala 94:53]
  assign Queue_108_clock = clock;
  assign Queue_108_reset = reset;
  assign Queue_108_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_44; // @[UserYanker.scala 95:53]
  assign Queue_108_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_108_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_108_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_44; // @[UserYanker.scala 94:53]
  assign Queue_109_clock = clock;
  assign Queue_109_reset = reset;
  assign Queue_109_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_45; // @[UserYanker.scala 95:53]
  assign Queue_109_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_109_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_109_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_45; // @[UserYanker.scala 94:53]
  assign Queue_110_clock = clock;
  assign Queue_110_reset = reset;
  assign Queue_110_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_46; // @[UserYanker.scala 95:53]
  assign Queue_110_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_110_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_110_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_46; // @[UserYanker.scala 94:53]
  assign Queue_111_clock = clock;
  assign Queue_111_reset = reset;
  assign Queue_111_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_47; // @[UserYanker.scala 95:53]
  assign Queue_111_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_111_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_111_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_47; // @[UserYanker.scala 94:53]
  assign Queue_112_clock = clock;
  assign Queue_112_reset = reset;
  assign Queue_112_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_48; // @[UserYanker.scala 95:53]
  assign Queue_112_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_112_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_112_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_48; // @[UserYanker.scala 94:53]
  assign Queue_113_clock = clock;
  assign Queue_113_reset = reset;
  assign Queue_113_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_49; // @[UserYanker.scala 95:53]
  assign Queue_113_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_113_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_113_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_49; // @[UserYanker.scala 94:53]
  assign Queue_114_clock = clock;
  assign Queue_114_reset = reset;
  assign Queue_114_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_50; // @[UserYanker.scala 95:53]
  assign Queue_114_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_114_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_114_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_50; // @[UserYanker.scala 94:53]
  assign Queue_115_clock = clock;
  assign Queue_115_reset = reset;
  assign Queue_115_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_51; // @[UserYanker.scala 95:53]
  assign Queue_115_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_115_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_115_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_51; // @[UserYanker.scala 94:53]
  assign Queue_116_clock = clock;
  assign Queue_116_reset = reset;
  assign Queue_116_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_52; // @[UserYanker.scala 95:53]
  assign Queue_116_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_116_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_116_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_52; // @[UserYanker.scala 94:53]
  assign Queue_117_clock = clock;
  assign Queue_117_reset = reset;
  assign Queue_117_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_53; // @[UserYanker.scala 95:53]
  assign Queue_117_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_117_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_117_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_53; // @[UserYanker.scala 94:53]
  assign Queue_118_clock = clock;
  assign Queue_118_reset = reset;
  assign Queue_118_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_54; // @[UserYanker.scala 95:53]
  assign Queue_118_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_118_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_118_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_54; // @[UserYanker.scala 94:53]
  assign Queue_119_clock = clock;
  assign Queue_119_reset = reset;
  assign Queue_119_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_55; // @[UserYanker.scala 95:53]
  assign Queue_119_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_119_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_119_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_55; // @[UserYanker.scala 94:53]
  assign Queue_120_clock = clock;
  assign Queue_120_reset = reset;
  assign Queue_120_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_56; // @[UserYanker.scala 95:53]
  assign Queue_120_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_120_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_120_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_56; // @[UserYanker.scala 94:53]
  assign Queue_121_clock = clock;
  assign Queue_121_reset = reset;
  assign Queue_121_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_57; // @[UserYanker.scala 95:53]
  assign Queue_121_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_121_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_121_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_57; // @[UserYanker.scala 94:53]
  assign Queue_122_clock = clock;
  assign Queue_122_reset = reset;
  assign Queue_122_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_58; // @[UserYanker.scala 95:53]
  assign Queue_122_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_122_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_122_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_58; // @[UserYanker.scala 94:53]
  assign Queue_123_clock = clock;
  assign Queue_123_reset = reset;
  assign Queue_123_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_59; // @[UserYanker.scala 95:53]
  assign Queue_123_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_123_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_123_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_59; // @[UserYanker.scala 94:53]
  assign Queue_124_clock = clock;
  assign Queue_124_reset = reset;
  assign Queue_124_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_60; // @[UserYanker.scala 95:53]
  assign Queue_124_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_124_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_124_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_60; // @[UserYanker.scala 94:53]
  assign Queue_125_clock = clock;
  assign Queue_125_reset = reset;
  assign Queue_125_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_61; // @[UserYanker.scala 95:53]
  assign Queue_125_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_125_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_125_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_61; // @[UserYanker.scala 94:53]
  assign Queue_126_clock = clock;
  assign Queue_126_reset = reset;
  assign Queue_126_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_62; // @[UserYanker.scala 95:53]
  assign Queue_126_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_126_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_126_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_62; // @[UserYanker.scala 94:53]
  assign Queue_127_clock = clock;
  assign Queue_127_reset = reset;
  assign Queue_127_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_63; // @[UserYanker.scala 95:53]
  assign Queue_127_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_127_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_127_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_63; // @[UserYanker.scala 94:53]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~auto_out_r_valid | _GEN_127)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at UserYanker.scala:66 assert (!out.r.valid || r_valid) // Q must be ready faster than the response\n"
            ); // @[UserYanker.scala 66:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~auto_out_r_valid | _GEN_127) & ~reset) begin
          $fatal; // @[UserYanker.scala 66:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3 & ~(~auto_out_b_valid | _GEN_447)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at UserYanker.scala:87 assert (!out.b.valid || b_valid) // Q must be ready faster than the response\n"
            ); // @[UserYanker.scala 87:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~auto_out_b_valid | _GEN_447) & _T_3) begin
          $fatal; // @[UserYanker.scala 87:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_161(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [5:0]  io_enq_bits_id,
  input  [33:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_len,
  input  [2:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_burst,
  input         io_enq_bits_lock,
  input  [3:0]  io_enq_bits_cache,
  input  [2:0]  io_enq_bits_prot,
  input  [3:0]  io_enq_bits_qos,
  input  [6:0]  io_enq_bits_echo_tl_state_source,
  input  [1:0]  io_enq_bits_echo_extra_id,
  input         io_deq_ready,
  output        io_deq_valid,
  output [5:0]  io_deq_bits_id,
  output [33:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_len,
  output [2:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_burst,
  output        io_deq_bits_lock,
  output [3:0]  io_deq_bits_cache,
  output [2:0]  io_deq_bits_prot,
  output [3:0]  io_deq_bits_qos,
  output [6:0]  io_deq_bits_echo_tl_state_source,
  output [1:0]  io_deq_bits_echo_extra_id
);
  reg [5:0] ram_id [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [5:0] ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [5:0] ram_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [33:0] ram_addr [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_addr_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_addr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [33:0] ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [33:0] ram_addr_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_addr_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_addr_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_addr_MPORT_en; // @[Decoupled.scala 273:95]
  reg [7:0] ram_len [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_len_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_len_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [7:0] ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [7:0] ram_len_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_len_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_len_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_len_MPORT_en; // @[Decoupled.scala 273:95]
  reg [2:0] ram_size [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_size_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_burst [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_burst_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_burst_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_burst_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_burst_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_burst_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_burst_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_lock [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_lock_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_lock_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_lock_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_lock_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_lock_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_lock_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_lock_MPORT_en; // @[Decoupled.scala 273:95]
  reg [3:0] ram_cache [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_cache_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_cache_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [3:0] ram_cache_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [3:0] ram_cache_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_cache_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_cache_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_cache_MPORT_en; // @[Decoupled.scala 273:95]
  reg [2:0] ram_prot [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_prot_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_prot_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [2:0] ram_prot_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_prot_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_prot_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_prot_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_prot_MPORT_en; // @[Decoupled.scala 273:95]
  reg [3:0] ram_qos [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_qos_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_qos_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [3:0] ram_qos_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [3:0] ram_qos_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_qos_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_qos_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_qos_MPORT_en; // @[Decoupled.scala 273:95]
  reg [6:0] ram_echo_tl_state_source [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [6:0] ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [6:0] ram_echo_tl_state_source_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_echo_extra_id [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_echo_extra_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_echo_extra_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_echo_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_echo_extra_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_echo_extra_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_echo_extra_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_echo_extra_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = enq_ptr_value;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_addr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_addr_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = enq_ptr_value;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_len_io_deq_bits_MPORT_en = 1'h1;
  assign ram_len_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_len_io_deq_bits_MPORT_data = ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_len_MPORT_data = io_enq_bits_len;
  assign ram_len_MPORT_addr = enq_ptr_value;
  assign ram_len_MPORT_mask = 1'h1;
  assign ram_len_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = enq_ptr_value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_burst_io_deq_bits_MPORT_en = 1'h1;
  assign ram_burst_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_burst_io_deq_bits_MPORT_data = ram_burst[ram_burst_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_burst_MPORT_data = io_enq_bits_burst;
  assign ram_burst_MPORT_addr = enq_ptr_value;
  assign ram_burst_MPORT_mask = 1'h1;
  assign ram_burst_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_lock_io_deq_bits_MPORT_en = 1'h1;
  assign ram_lock_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_lock_io_deq_bits_MPORT_data = ram_lock[ram_lock_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_lock_MPORT_data = io_enq_bits_lock;
  assign ram_lock_MPORT_addr = enq_ptr_value;
  assign ram_lock_MPORT_mask = 1'h1;
  assign ram_lock_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_cache_io_deq_bits_MPORT_en = 1'h1;
  assign ram_cache_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_cache_io_deq_bits_MPORT_data = ram_cache[ram_cache_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_cache_MPORT_data = io_enq_bits_cache;
  assign ram_cache_MPORT_addr = enq_ptr_value;
  assign ram_cache_MPORT_mask = 1'h1;
  assign ram_cache_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_prot_io_deq_bits_MPORT_en = 1'h1;
  assign ram_prot_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_prot_io_deq_bits_MPORT_data = ram_prot[ram_prot_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_prot_MPORT_data = io_enq_bits_prot;
  assign ram_prot_MPORT_addr = enq_ptr_value;
  assign ram_prot_MPORT_mask = 1'h1;
  assign ram_prot_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_qos_io_deq_bits_MPORT_en = 1'h1;
  assign ram_qos_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_qos_io_deq_bits_MPORT_data = ram_qos[ram_qos_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_qos_MPORT_data = io_enq_bits_qos;
  assign ram_qos_MPORT_addr = enq_ptr_value;
  assign ram_qos_MPORT_mask = 1'h1;
  assign ram_qos_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_data =
    ram_echo_tl_state_source[ram_echo_tl_state_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_echo_tl_state_source_MPORT_data = io_enq_bits_echo_tl_state_source;
  assign ram_echo_tl_state_source_MPORT_addr = enq_ptr_value;
  assign ram_echo_tl_state_source_MPORT_mask = 1'h1;
  assign ram_echo_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_echo_extra_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_echo_extra_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_echo_extra_id_io_deq_bits_MPORT_data = ram_echo_extra_id[ram_echo_extra_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_echo_extra_id_MPORT_data = io_enq_bits_echo_extra_id;
  assign ram_echo_extra_id_MPORT_addr = enq_ptr_value;
  assign ram_echo_extra_id_MPORT_mask = 1'h1;
  assign ram_echo_extra_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_id = ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_addr = ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_len = ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_burst = ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_lock = ram_lock_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_cache = ram_cache_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_prot = ram_prot_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_qos = ram_qos_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_echo_tl_state_source = ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_echo_extra_id = ram_echo_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_len_MPORT_en & ram_len_MPORT_mask) begin
      ram_len[ram_len_MPORT_addr] <= ram_len_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_burst_MPORT_en & ram_burst_MPORT_mask) begin
      ram_burst[ram_burst_MPORT_addr] <= ram_burst_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_lock_MPORT_en & ram_lock_MPORT_mask) begin
      ram_lock[ram_lock_MPORT_addr] <= ram_lock_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_cache_MPORT_en & ram_cache_MPORT_mask) begin
      ram_cache[ram_cache_MPORT_addr] <= ram_cache_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_prot_MPORT_en & ram_prot_MPORT_mask) begin
      ram_prot[ram_prot_MPORT_addr] <= ram_prot_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_qos_MPORT_en & ram_qos_MPORT_mask) begin
      ram_qos[ram_qos_MPORT_addr] <= ram_qos_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_echo_tl_state_source_MPORT_en & ram_echo_tl_state_source_MPORT_mask) begin
      ram_echo_tl_state_source[ram_echo_tl_state_source_MPORT_addr] <= ram_echo_tl_state_source_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_echo_extra_id_MPORT_en & ram_echo_extra_id_MPORT_mask) begin
      ram_echo_extra_id[ram_echo_extra_id_MPORT_addr] <= ram_echo_extra_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
endmodule
module Queue_163(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [5:0] io_enq_bits_id,
  input  [1:0] io_enq_bits_resp,
  input  [6:0] io_enq_bits_echo_tl_state_source,
  input  [1:0] io_enq_bits_echo_extra_id,
  input        io_deq_ready,
  output       io_deq_valid,
  output [5:0] io_deq_bits_id,
  output [1:0] io_deq_bits_resp,
  output [6:0] io_deq_bits_echo_tl_state_source,
  output [1:0] io_deq_bits_echo_extra_id
);
  reg [5:0] ram_id [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [5:0] ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [5:0] ram_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_resp [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_resp_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_resp_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_resp_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_en; // @[Decoupled.scala 273:95]
  reg [6:0] ram_echo_tl_state_source [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [6:0] ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [6:0] ram_echo_tl_state_source_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_echo_extra_id [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_echo_extra_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_echo_extra_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_echo_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_echo_extra_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_echo_extra_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_echo_extra_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_echo_extra_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = enq_ptr_value;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_resp_io_deq_bits_MPORT_en = 1'h1;
  assign ram_resp_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_resp_io_deq_bits_MPORT_data = ram_resp[ram_resp_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_resp_MPORT_data = io_enq_bits_resp;
  assign ram_resp_MPORT_addr = enq_ptr_value;
  assign ram_resp_MPORT_mask = 1'h1;
  assign ram_resp_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_data =
    ram_echo_tl_state_source[ram_echo_tl_state_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_echo_tl_state_source_MPORT_data = io_enq_bits_echo_tl_state_source;
  assign ram_echo_tl_state_source_MPORT_addr = enq_ptr_value;
  assign ram_echo_tl_state_source_MPORT_mask = 1'h1;
  assign ram_echo_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_echo_extra_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_echo_extra_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_echo_extra_id_io_deq_bits_MPORT_data = ram_echo_extra_id[ram_echo_extra_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_echo_extra_id_MPORT_data = io_enq_bits_echo_extra_id;
  assign ram_echo_extra_id_MPORT_addr = enq_ptr_value;
  assign ram_echo_extra_id_MPORT_mask = 1'h1;
  assign ram_echo_extra_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_id = ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_resp = ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_echo_tl_state_source = ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_echo_extra_id = ram_echo_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_resp_MPORT_en & ram_resp_MPORT_mask) begin
      ram_resp[ram_resp_MPORT_addr] <= ram_resp_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_echo_tl_state_source_MPORT_en & ram_echo_tl_state_source_MPORT_mask) begin
      ram_echo_tl_state_source[ram_echo_tl_state_source_MPORT_addr] <= ram_echo_tl_state_source_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_echo_extra_id_MPORT_en & ram_echo_extra_id_MPORT_mask) begin
      ram_echo_extra_id[ram_echo_extra_id_MPORT_addr] <= ram_echo_extra_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
endmodule
module Queue_165(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [5:0]   io_enq_bits_id,
  input  [511:0] io_enq_bits_data,
  input  [1:0]   io_enq_bits_resp,
  input  [6:0]   io_enq_bits_echo_tl_state_source,
  input  [1:0]   io_enq_bits_echo_extra_id,
  input          io_enq_bits_last,
  input          io_deq_ready,
  output         io_deq_valid,
  output [5:0]   io_deq_bits_id,
  output [511:0] io_deq_bits_data,
  output [1:0]   io_deq_bits_resp,
  output [6:0]   io_deq_bits_echo_tl_state_source,
  output [1:0]   io_deq_bits_echo_extra_id,
  output         io_deq_bits_last
);
  reg [5:0] ram_id [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [5:0] ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [5:0] ram_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [511:0] ram_data [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [511:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [511:0] ram_data_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_resp [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_resp_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_resp_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_resp_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_en; // @[Decoupled.scala 273:95]
  reg [6:0] ram_echo_tl_state_source [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [6:0] ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [6:0] ram_echo_tl_state_source_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_echo_extra_id [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_echo_extra_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_echo_extra_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_echo_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_echo_extra_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_echo_extra_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_echo_extra_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_echo_extra_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_last [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = enq_ptr_value;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_resp_io_deq_bits_MPORT_en = 1'h1;
  assign ram_resp_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_resp_io_deq_bits_MPORT_data = ram_resp[ram_resp_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_resp_MPORT_data = io_enq_bits_resp;
  assign ram_resp_MPORT_addr = enq_ptr_value;
  assign ram_resp_MPORT_mask = 1'h1;
  assign ram_resp_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_data =
    ram_echo_tl_state_source[ram_echo_tl_state_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_echo_tl_state_source_MPORT_data = io_enq_bits_echo_tl_state_source;
  assign ram_echo_tl_state_source_MPORT_addr = enq_ptr_value;
  assign ram_echo_tl_state_source_MPORT_mask = 1'h1;
  assign ram_echo_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_echo_extra_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_echo_extra_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_echo_extra_id_io_deq_bits_MPORT_data = ram_echo_extra_id[ram_echo_extra_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_echo_extra_id_MPORT_data = io_enq_bits_echo_extra_id;
  assign ram_echo_extra_id_MPORT_addr = enq_ptr_value;
  assign ram_echo_extra_id_MPORT_mask = 1'h1;
  assign ram_echo_extra_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_last_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_last_io_deq_bits_MPORT_data = ram_last[ram_last_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_last_MPORT_data = io_enq_bits_last;
  assign ram_last_MPORT_addr = enq_ptr_value;
  assign ram_last_MPORT_mask = 1'h1;
  assign ram_last_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_id = ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_resp = ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_echo_tl_state_source = ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_echo_extra_id = ram_echo_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_last = ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_resp_MPORT_en & ram_resp_MPORT_mask) begin
      ram_resp[ram_resp_MPORT_addr] <= ram_resp_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_echo_tl_state_source_MPORT_en & ram_echo_tl_state_source_MPORT_mask) begin
      ram_echo_tl_state_source[ram_echo_tl_state_source_MPORT_addr] <= ram_echo_tl_state_source_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_echo_extra_id_MPORT_en & ram_echo_extra_id_MPORT_mask) begin
      ram_echo_extra_id[ram_echo_extra_id_MPORT_addr] <= ram_echo_extra_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_last_MPORT_en & ram_last_MPORT_mask) begin
      ram_last[ram_last_MPORT_addr] <= ram_last_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
endmodule
module AXI4Buffer_4(
  input          clock,
  input          reset,
  output         auto_in_aw_ready,
  input          auto_in_aw_valid,
  input  [5:0]   auto_in_aw_bits_id,
  input  [33:0]  auto_in_aw_bits_addr,
  input  [7:0]   auto_in_aw_bits_len,
  input  [2:0]   auto_in_aw_bits_size,
  input  [1:0]   auto_in_aw_bits_burst,
  input          auto_in_aw_bits_lock,
  input  [3:0]   auto_in_aw_bits_cache,
  input  [2:0]   auto_in_aw_bits_prot,
  input  [3:0]   auto_in_aw_bits_qos,
  input  [6:0]   auto_in_aw_bits_echo_tl_state_source,
  input  [1:0]   auto_in_aw_bits_echo_extra_id,
  output         auto_in_w_ready,
  input          auto_in_w_valid,
  input  [511:0] auto_in_w_bits_data,
  input  [63:0]  auto_in_w_bits_strb,
  input          auto_in_w_bits_last,
  input          auto_in_b_ready,
  output         auto_in_b_valid,
  output [5:0]   auto_in_b_bits_id,
  output [1:0]   auto_in_b_bits_resp,
  output [6:0]   auto_in_b_bits_echo_tl_state_source,
  output [1:0]   auto_in_b_bits_echo_extra_id,
  output         auto_in_ar_ready,
  input          auto_in_ar_valid,
  input  [5:0]   auto_in_ar_bits_id,
  input  [33:0]  auto_in_ar_bits_addr,
  input  [7:0]   auto_in_ar_bits_len,
  input  [2:0]   auto_in_ar_bits_size,
  input  [1:0]   auto_in_ar_bits_burst,
  input          auto_in_ar_bits_lock,
  input  [3:0]   auto_in_ar_bits_cache,
  input  [2:0]   auto_in_ar_bits_prot,
  input  [3:0]   auto_in_ar_bits_qos,
  input  [6:0]   auto_in_ar_bits_echo_tl_state_source,
  input  [1:0]   auto_in_ar_bits_echo_extra_id,
  input          auto_in_r_ready,
  output         auto_in_r_valid,
  output [5:0]   auto_in_r_bits_id,
  output [511:0] auto_in_r_bits_data,
  output [1:0]   auto_in_r_bits_resp,
  output [6:0]   auto_in_r_bits_echo_tl_state_source,
  output [1:0]   auto_in_r_bits_echo_extra_id,
  output         auto_in_r_bits_last,
  input          auto_out_aw_ready,
  output         auto_out_aw_valid,
  output [5:0]   auto_out_aw_bits_id,
  output [33:0]  auto_out_aw_bits_addr,
  output [7:0]   auto_out_aw_bits_len,
  output [2:0]   auto_out_aw_bits_size,
  output [1:0]   auto_out_aw_bits_burst,
  output         auto_out_aw_bits_lock,
  output [3:0]   auto_out_aw_bits_cache,
  output [2:0]   auto_out_aw_bits_prot,
  output [3:0]   auto_out_aw_bits_qos,
  output [6:0]   auto_out_aw_bits_echo_tl_state_source,
  output [1:0]   auto_out_aw_bits_echo_extra_id,
  input          auto_out_w_ready,
  output         auto_out_w_valid,
  output [511:0] auto_out_w_bits_data,
  output [63:0]  auto_out_w_bits_strb,
  output         auto_out_w_bits_last,
  output         auto_out_b_ready,
  input          auto_out_b_valid,
  input  [5:0]   auto_out_b_bits_id,
  input  [1:0]   auto_out_b_bits_resp,
  input  [6:0]   auto_out_b_bits_echo_tl_state_source,
  input  [1:0]   auto_out_b_bits_echo_extra_id,
  input          auto_out_ar_ready,
  output         auto_out_ar_valid,
  output [5:0]   auto_out_ar_bits_id,
  output [33:0]  auto_out_ar_bits_addr,
  output [7:0]   auto_out_ar_bits_len,
  output [2:0]   auto_out_ar_bits_size,
  output [1:0]   auto_out_ar_bits_burst,
  output         auto_out_ar_bits_lock,
  output [3:0]   auto_out_ar_bits_cache,
  output [2:0]   auto_out_ar_bits_prot,
  output [3:0]   auto_out_ar_bits_qos,
  output [6:0]   auto_out_ar_bits_echo_tl_state_source,
  output [1:0]   auto_out_ar_bits_echo_extra_id,
  output         auto_out_r_ready,
  input          auto_out_r_valid,
  input  [5:0]   auto_out_r_bits_id,
  input  [511:0] auto_out_r_bits_data,
  input  [1:0]   auto_out_r_bits_resp,
  input  [6:0]   auto_out_r_bits_echo_tl_state_source,
  input  [1:0]   auto_out_r_bits_echo_extra_id,
  input          auto_out_r_bits_last
);
  wire  x1_aw_deq_clock; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_reset; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [5:0] x1_aw_deq_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire [33:0] x1_aw_deq_io_enq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] x1_aw_deq_io_enq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] x1_aw_deq_io_enq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] x1_aw_deq_io_enq_bits_burst; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_enq_bits_lock; // @[Decoupled.scala 375:21]
  wire [3:0] x1_aw_deq_io_enq_bits_cache; // @[Decoupled.scala 375:21]
  wire [2:0] x1_aw_deq_io_enq_bits_prot; // @[Decoupled.scala 375:21]
  wire [3:0] x1_aw_deq_io_enq_bits_qos; // @[Decoupled.scala 375:21]
  wire [6:0] x1_aw_deq_io_enq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire [1:0] x1_aw_deq_io_enq_bits_echo_extra_id; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [5:0] x1_aw_deq_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [33:0] x1_aw_deq_io_deq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] x1_aw_deq_io_deq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] x1_aw_deq_io_deq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] x1_aw_deq_io_deq_bits_burst; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_deq_bits_lock; // @[Decoupled.scala 375:21]
  wire [3:0] x1_aw_deq_io_deq_bits_cache; // @[Decoupled.scala 375:21]
  wire [2:0] x1_aw_deq_io_deq_bits_prot; // @[Decoupled.scala 375:21]
  wire [3:0] x1_aw_deq_io_deq_bits_qos; // @[Decoupled.scala 375:21]
  wire [6:0] x1_aw_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire [1:0] x1_aw_deq_io_deq_bits_echo_extra_id; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_clock; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_reset; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [511:0] x1_w_deq_io_enq_bits_data; // @[Decoupled.scala 375:21]
  wire [63:0] x1_w_deq_io_enq_bits_strb; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_enq_bits_last; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [511:0] x1_w_deq_io_deq_bits_data; // @[Decoupled.scala 375:21]
  wire [63:0] x1_w_deq_io_deq_bits_strb; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_deq_bits_last; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_clock; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_reset; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [5:0] bundleIn_0_b_deq_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire [1:0] bundleIn_0_b_deq_io_enq_bits_resp; // @[Decoupled.scala 375:21]
  wire [6:0] bundleIn_0_b_deq_io_enq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire [1:0] bundleIn_0_b_deq_io_enq_bits_echo_extra_id; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [5:0] bundleIn_0_b_deq_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [1:0] bundleIn_0_b_deq_io_deq_bits_resp; // @[Decoupled.scala 375:21]
  wire [6:0] bundleIn_0_b_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire [1:0] bundleIn_0_b_deq_io_deq_bits_echo_extra_id; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_clock; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_reset; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [5:0] x1_ar_deq_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire [33:0] x1_ar_deq_io_enq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] x1_ar_deq_io_enq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] x1_ar_deq_io_enq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] x1_ar_deq_io_enq_bits_burst; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_enq_bits_lock; // @[Decoupled.scala 375:21]
  wire [3:0] x1_ar_deq_io_enq_bits_cache; // @[Decoupled.scala 375:21]
  wire [2:0] x1_ar_deq_io_enq_bits_prot; // @[Decoupled.scala 375:21]
  wire [3:0] x1_ar_deq_io_enq_bits_qos; // @[Decoupled.scala 375:21]
  wire [6:0] x1_ar_deq_io_enq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire [1:0] x1_ar_deq_io_enq_bits_echo_extra_id; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [5:0] x1_ar_deq_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [33:0] x1_ar_deq_io_deq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] x1_ar_deq_io_deq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] x1_ar_deq_io_deq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] x1_ar_deq_io_deq_bits_burst; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_deq_bits_lock; // @[Decoupled.scala 375:21]
  wire [3:0] x1_ar_deq_io_deq_bits_cache; // @[Decoupled.scala 375:21]
  wire [2:0] x1_ar_deq_io_deq_bits_prot; // @[Decoupled.scala 375:21]
  wire [3:0] x1_ar_deq_io_deq_bits_qos; // @[Decoupled.scala 375:21]
  wire [6:0] x1_ar_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire [1:0] x1_ar_deq_io_deq_bits_echo_extra_id; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_clock; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_reset; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [5:0] bundleIn_0_r_deq_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire [511:0] bundleIn_0_r_deq_io_enq_bits_data; // @[Decoupled.scala 375:21]
  wire [1:0] bundleIn_0_r_deq_io_enq_bits_resp; // @[Decoupled.scala 375:21]
  wire [6:0] bundleIn_0_r_deq_io_enq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire [1:0] bundleIn_0_r_deq_io_enq_bits_echo_extra_id; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_enq_bits_last; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [5:0] bundleIn_0_r_deq_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [511:0] bundleIn_0_r_deq_io_deq_bits_data; // @[Decoupled.scala 375:21]
  wire [1:0] bundleIn_0_r_deq_io_deq_bits_resp; // @[Decoupled.scala 375:21]
  wire [6:0] bundleIn_0_r_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire [1:0] bundleIn_0_r_deq_io_deq_bits_echo_extra_id; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_deq_bits_last; // @[Decoupled.scala 375:21]
  Queue_161 x1_aw_deq ( // @[Decoupled.scala 375:21]
    .clock(x1_aw_deq_clock),
    .reset(x1_aw_deq_reset),
    .io_enq_ready(x1_aw_deq_io_enq_ready),
    .io_enq_valid(x1_aw_deq_io_enq_valid),
    .io_enq_bits_id(x1_aw_deq_io_enq_bits_id),
    .io_enq_bits_addr(x1_aw_deq_io_enq_bits_addr),
    .io_enq_bits_len(x1_aw_deq_io_enq_bits_len),
    .io_enq_bits_size(x1_aw_deq_io_enq_bits_size),
    .io_enq_bits_burst(x1_aw_deq_io_enq_bits_burst),
    .io_enq_bits_lock(x1_aw_deq_io_enq_bits_lock),
    .io_enq_bits_cache(x1_aw_deq_io_enq_bits_cache),
    .io_enq_bits_prot(x1_aw_deq_io_enq_bits_prot),
    .io_enq_bits_qos(x1_aw_deq_io_enq_bits_qos),
    .io_enq_bits_echo_tl_state_source(x1_aw_deq_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_echo_extra_id(x1_aw_deq_io_enq_bits_echo_extra_id),
    .io_deq_ready(x1_aw_deq_io_deq_ready),
    .io_deq_valid(x1_aw_deq_io_deq_valid),
    .io_deq_bits_id(x1_aw_deq_io_deq_bits_id),
    .io_deq_bits_addr(x1_aw_deq_io_deq_bits_addr),
    .io_deq_bits_len(x1_aw_deq_io_deq_bits_len),
    .io_deq_bits_size(x1_aw_deq_io_deq_bits_size),
    .io_deq_bits_burst(x1_aw_deq_io_deq_bits_burst),
    .io_deq_bits_lock(x1_aw_deq_io_deq_bits_lock),
    .io_deq_bits_cache(x1_aw_deq_io_deq_bits_cache),
    .io_deq_bits_prot(x1_aw_deq_io_deq_bits_prot),
    .io_deq_bits_qos(x1_aw_deq_io_deq_bits_qos),
    .io_deq_bits_echo_tl_state_source(x1_aw_deq_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_echo_extra_id(x1_aw_deq_io_deq_bits_echo_extra_id)
  );
  Queue_7 x1_w_deq ( // @[Decoupled.scala 375:21]
    .clock(x1_w_deq_clock),
    .reset(x1_w_deq_reset),
    .io_enq_ready(x1_w_deq_io_enq_ready),
    .io_enq_valid(x1_w_deq_io_enq_valid),
    .io_enq_bits_data(x1_w_deq_io_enq_bits_data),
    .io_enq_bits_strb(x1_w_deq_io_enq_bits_strb),
    .io_enq_bits_last(x1_w_deq_io_enq_bits_last),
    .io_deq_ready(x1_w_deq_io_deq_ready),
    .io_deq_valid(x1_w_deq_io_deq_valid),
    .io_deq_bits_data(x1_w_deq_io_deq_bits_data),
    .io_deq_bits_strb(x1_w_deq_io_deq_bits_strb),
    .io_deq_bits_last(x1_w_deq_io_deq_bits_last)
  );
  Queue_163 bundleIn_0_b_deq ( // @[Decoupled.scala 375:21]
    .clock(bundleIn_0_b_deq_clock),
    .reset(bundleIn_0_b_deq_reset),
    .io_enq_ready(bundleIn_0_b_deq_io_enq_ready),
    .io_enq_valid(bundleIn_0_b_deq_io_enq_valid),
    .io_enq_bits_id(bundleIn_0_b_deq_io_enq_bits_id),
    .io_enq_bits_resp(bundleIn_0_b_deq_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_source(bundleIn_0_b_deq_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_echo_extra_id(bundleIn_0_b_deq_io_enq_bits_echo_extra_id),
    .io_deq_ready(bundleIn_0_b_deq_io_deq_ready),
    .io_deq_valid(bundleIn_0_b_deq_io_deq_valid),
    .io_deq_bits_id(bundleIn_0_b_deq_io_deq_bits_id),
    .io_deq_bits_resp(bundleIn_0_b_deq_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_source(bundleIn_0_b_deq_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_echo_extra_id(bundleIn_0_b_deq_io_deq_bits_echo_extra_id)
  );
  Queue_161 x1_ar_deq ( // @[Decoupled.scala 375:21]
    .clock(x1_ar_deq_clock),
    .reset(x1_ar_deq_reset),
    .io_enq_ready(x1_ar_deq_io_enq_ready),
    .io_enq_valid(x1_ar_deq_io_enq_valid),
    .io_enq_bits_id(x1_ar_deq_io_enq_bits_id),
    .io_enq_bits_addr(x1_ar_deq_io_enq_bits_addr),
    .io_enq_bits_len(x1_ar_deq_io_enq_bits_len),
    .io_enq_bits_size(x1_ar_deq_io_enq_bits_size),
    .io_enq_bits_burst(x1_ar_deq_io_enq_bits_burst),
    .io_enq_bits_lock(x1_ar_deq_io_enq_bits_lock),
    .io_enq_bits_cache(x1_ar_deq_io_enq_bits_cache),
    .io_enq_bits_prot(x1_ar_deq_io_enq_bits_prot),
    .io_enq_bits_qos(x1_ar_deq_io_enq_bits_qos),
    .io_enq_bits_echo_tl_state_source(x1_ar_deq_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_echo_extra_id(x1_ar_deq_io_enq_bits_echo_extra_id),
    .io_deq_ready(x1_ar_deq_io_deq_ready),
    .io_deq_valid(x1_ar_deq_io_deq_valid),
    .io_deq_bits_id(x1_ar_deq_io_deq_bits_id),
    .io_deq_bits_addr(x1_ar_deq_io_deq_bits_addr),
    .io_deq_bits_len(x1_ar_deq_io_deq_bits_len),
    .io_deq_bits_size(x1_ar_deq_io_deq_bits_size),
    .io_deq_bits_burst(x1_ar_deq_io_deq_bits_burst),
    .io_deq_bits_lock(x1_ar_deq_io_deq_bits_lock),
    .io_deq_bits_cache(x1_ar_deq_io_deq_bits_cache),
    .io_deq_bits_prot(x1_ar_deq_io_deq_bits_prot),
    .io_deq_bits_qos(x1_ar_deq_io_deq_bits_qos),
    .io_deq_bits_echo_tl_state_source(x1_ar_deq_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_echo_extra_id(x1_ar_deq_io_deq_bits_echo_extra_id)
  );
  Queue_165 bundleIn_0_r_deq ( // @[Decoupled.scala 375:21]
    .clock(bundleIn_0_r_deq_clock),
    .reset(bundleIn_0_r_deq_reset),
    .io_enq_ready(bundleIn_0_r_deq_io_enq_ready),
    .io_enq_valid(bundleIn_0_r_deq_io_enq_valid),
    .io_enq_bits_id(bundleIn_0_r_deq_io_enq_bits_id),
    .io_enq_bits_data(bundleIn_0_r_deq_io_enq_bits_data),
    .io_enq_bits_resp(bundleIn_0_r_deq_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_source(bundleIn_0_r_deq_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_echo_extra_id(bundleIn_0_r_deq_io_enq_bits_echo_extra_id),
    .io_enq_bits_last(bundleIn_0_r_deq_io_enq_bits_last),
    .io_deq_ready(bundleIn_0_r_deq_io_deq_ready),
    .io_deq_valid(bundleIn_0_r_deq_io_deq_valid),
    .io_deq_bits_id(bundleIn_0_r_deq_io_deq_bits_id),
    .io_deq_bits_data(bundleIn_0_r_deq_io_deq_bits_data),
    .io_deq_bits_resp(bundleIn_0_r_deq_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_source(bundleIn_0_r_deq_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_echo_extra_id(bundleIn_0_r_deq_io_deq_bits_echo_extra_id),
    .io_deq_bits_last(bundleIn_0_r_deq_io_deq_bits_last)
  );
  assign auto_in_aw_ready = x1_aw_deq_io_enq_ready; // @[Nodes.scala 1215:84 Decoupled.scala 379:17]
  assign auto_in_w_ready = x1_w_deq_io_enq_ready; // @[Nodes.scala 1215:84 Decoupled.scala 379:17]
  assign auto_in_b_valid = bundleIn_0_b_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_in_b_bits_id = bundleIn_0_b_deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_b_bits_resp = bundleIn_0_b_deq_io_deq_bits_resp; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_b_bits_echo_tl_state_source = bundleIn_0_b_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_b_bits_echo_extra_id = bundleIn_0_b_deq_io_deq_bits_echo_extra_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_ar_ready = x1_ar_deq_io_enq_ready; // @[Nodes.scala 1215:84 Decoupled.scala 379:17]
  assign auto_in_r_valid = bundleIn_0_r_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_in_r_bits_id = bundleIn_0_r_deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_r_bits_data = bundleIn_0_r_deq_io_deq_bits_data; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_r_bits_resp = bundleIn_0_r_deq_io_deq_bits_resp; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_r_bits_echo_tl_state_source = bundleIn_0_r_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_r_bits_echo_extra_id = bundleIn_0_r_deq_io_deq_bits_echo_extra_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_r_bits_last = bundleIn_0_r_deq_io_deq_bits_last; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_valid = x1_aw_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_out_aw_bits_id = x1_aw_deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_addr = x1_aw_deq_io_deq_bits_addr; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_len = x1_aw_deq_io_deq_bits_len; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_size = x1_aw_deq_io_deq_bits_size; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_burst = x1_aw_deq_io_deq_bits_burst; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_lock = x1_aw_deq_io_deq_bits_lock; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_cache = x1_aw_deq_io_deq_bits_cache; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_prot = x1_aw_deq_io_deq_bits_prot; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_qos = x1_aw_deq_io_deq_bits_qos; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_echo_tl_state_source = x1_aw_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_echo_extra_id = x1_aw_deq_io_deq_bits_echo_extra_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_w_valid = x1_w_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_out_w_bits_data = x1_w_deq_io_deq_bits_data; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_w_bits_strb = x1_w_deq_io_deq_bits_strb; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_w_bits_last = x1_w_deq_io_deq_bits_last; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_b_ready = bundleIn_0_b_deq_io_enq_ready; // @[Nodes.scala 1212:84 Decoupled.scala 379:17]
  assign auto_out_ar_valid = x1_ar_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_out_ar_bits_id = x1_ar_deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_addr = x1_ar_deq_io_deq_bits_addr; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_len = x1_ar_deq_io_deq_bits_len; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_size = x1_ar_deq_io_deq_bits_size; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_burst = x1_ar_deq_io_deq_bits_burst; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_lock = x1_ar_deq_io_deq_bits_lock; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_cache = x1_ar_deq_io_deq_bits_cache; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_prot = x1_ar_deq_io_deq_bits_prot; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_qos = x1_ar_deq_io_deq_bits_qos; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_echo_tl_state_source = x1_ar_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_echo_extra_id = x1_ar_deq_io_deq_bits_echo_extra_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_r_ready = bundleIn_0_r_deq_io_enq_ready; // @[Nodes.scala 1212:84 Decoupled.scala 379:17]
  assign x1_aw_deq_clock = clock;
  assign x1_aw_deq_reset = reset;
  assign x1_aw_deq_io_enq_valid = auto_in_aw_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_id = auto_in_aw_bits_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_addr = auto_in_aw_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_len = auto_in_aw_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_size = auto_in_aw_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_burst = auto_in_aw_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_lock = auto_in_aw_bits_lock; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_cache = auto_in_aw_bits_cache; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_prot = auto_in_aw_bits_prot; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_qos = auto_in_aw_bits_qos; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_echo_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_echo_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_deq_ready = auto_out_aw_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign x1_w_deq_clock = clock;
  assign x1_w_deq_reset = reset;
  assign x1_w_deq_io_enq_valid = auto_in_w_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_w_deq_io_enq_bits_data = auto_in_w_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_w_deq_io_enq_bits_strb = auto_in_w_bits_strb; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_w_deq_io_enq_bits_last = auto_in_w_bits_last; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_w_deq_io_deq_ready = auto_out_w_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_b_deq_clock = clock;
  assign bundleIn_0_b_deq_reset = reset;
  assign bundleIn_0_b_deq_io_enq_valid = auto_out_b_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_b_deq_io_enq_bits_id = auto_out_b_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_b_deq_io_enq_bits_resp = auto_out_b_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_b_deq_io_enq_bits_echo_tl_state_source = auto_out_b_bits_echo_tl_state_source; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_b_deq_io_enq_bits_echo_extra_id = auto_out_b_bits_echo_extra_id; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_b_deq_io_deq_ready = auto_in_b_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_clock = clock;
  assign x1_ar_deq_reset = reset;
  assign x1_ar_deq_io_enq_valid = auto_in_ar_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_id = auto_in_ar_bits_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_addr = auto_in_ar_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_len = auto_in_ar_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_size = auto_in_ar_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_burst = auto_in_ar_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_lock = auto_in_ar_bits_lock; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_cache = auto_in_ar_bits_cache; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_prot = auto_in_ar_bits_prot; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_qos = auto_in_ar_bits_qos; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_echo_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_echo_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_deq_ready = auto_out_ar_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_clock = clock;
  assign bundleIn_0_r_deq_reset = reset;
  assign bundleIn_0_r_deq_io_enq_valid = auto_out_r_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_enq_bits_id = auto_out_r_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_enq_bits_data = auto_out_r_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_enq_bits_resp = auto_out_r_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_enq_bits_echo_tl_state_source = auto_out_r_bits_echo_tl_state_source; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_enq_bits_echo_extra_id = auto_out_r_bits_echo_extra_id; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_enq_bits_last = auto_out_r_bits_last; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_deq_ready = auto_in_r_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
endmodule
module AXI4IdIndexer(
  output         auto_in_aw_ready,
  input          auto_in_aw_valid,
  input  [7:0]   auto_in_aw_bits_id,
  input  [33:0]  auto_in_aw_bits_addr,
  input  [7:0]   auto_in_aw_bits_len,
  input  [2:0]   auto_in_aw_bits_size,
  input  [1:0]   auto_in_aw_bits_burst,
  input          auto_in_aw_bits_lock,
  input  [3:0]   auto_in_aw_bits_cache,
  input  [2:0]   auto_in_aw_bits_prot,
  input  [3:0]   auto_in_aw_bits_qos,
  input  [6:0]   auto_in_aw_bits_echo_tl_state_source,
  output         auto_in_w_ready,
  input          auto_in_w_valid,
  input  [511:0] auto_in_w_bits_data,
  input  [63:0]  auto_in_w_bits_strb,
  input          auto_in_w_bits_last,
  input          auto_in_b_ready,
  output         auto_in_b_valid,
  output [7:0]   auto_in_b_bits_id,
  output [1:0]   auto_in_b_bits_resp,
  output [6:0]   auto_in_b_bits_echo_tl_state_source,
  output         auto_in_ar_ready,
  input          auto_in_ar_valid,
  input  [7:0]   auto_in_ar_bits_id,
  input  [33:0]  auto_in_ar_bits_addr,
  input  [7:0]   auto_in_ar_bits_len,
  input  [2:0]   auto_in_ar_bits_size,
  input  [1:0]   auto_in_ar_bits_burst,
  input          auto_in_ar_bits_lock,
  input  [3:0]   auto_in_ar_bits_cache,
  input  [2:0]   auto_in_ar_bits_prot,
  input  [3:0]   auto_in_ar_bits_qos,
  input  [6:0]   auto_in_ar_bits_echo_tl_state_source,
  input          auto_in_r_ready,
  output         auto_in_r_valid,
  output [7:0]   auto_in_r_bits_id,
  output [511:0] auto_in_r_bits_data,
  output [1:0]   auto_in_r_bits_resp,
  output [6:0]   auto_in_r_bits_echo_tl_state_source,
  output         auto_in_r_bits_last,
  input          auto_out_aw_ready,
  output         auto_out_aw_valid,
  output [5:0]   auto_out_aw_bits_id,
  output [33:0]  auto_out_aw_bits_addr,
  output [7:0]   auto_out_aw_bits_len,
  output [2:0]   auto_out_aw_bits_size,
  output [1:0]   auto_out_aw_bits_burst,
  output         auto_out_aw_bits_lock,
  output [3:0]   auto_out_aw_bits_cache,
  output [2:0]   auto_out_aw_bits_prot,
  output [3:0]   auto_out_aw_bits_qos,
  output [6:0]   auto_out_aw_bits_echo_tl_state_source,
  output [1:0]   auto_out_aw_bits_echo_extra_id,
  input          auto_out_w_ready,
  output         auto_out_w_valid,
  output [511:0] auto_out_w_bits_data,
  output [63:0]  auto_out_w_bits_strb,
  output         auto_out_w_bits_last,
  output         auto_out_b_ready,
  input          auto_out_b_valid,
  input  [5:0]   auto_out_b_bits_id,
  input  [1:0]   auto_out_b_bits_resp,
  input  [6:0]   auto_out_b_bits_echo_tl_state_source,
  input  [1:0]   auto_out_b_bits_echo_extra_id,
  input          auto_out_ar_ready,
  output         auto_out_ar_valid,
  output [5:0]   auto_out_ar_bits_id,
  output [33:0]  auto_out_ar_bits_addr,
  output [7:0]   auto_out_ar_bits_len,
  output [2:0]   auto_out_ar_bits_size,
  output [1:0]   auto_out_ar_bits_burst,
  output         auto_out_ar_bits_lock,
  output [3:0]   auto_out_ar_bits_cache,
  output [2:0]   auto_out_ar_bits_prot,
  output [3:0]   auto_out_ar_bits_qos,
  output [6:0]   auto_out_ar_bits_echo_tl_state_source,
  output [1:0]   auto_out_ar_bits_echo_extra_id,
  output         auto_out_r_ready,
  input          auto_out_r_valid,
  input  [5:0]   auto_out_r_bits_id,
  input  [511:0] auto_out_r_bits_data,
  input  [1:0]   auto_out_r_bits_resp,
  input  [6:0]   auto_out_r_bits_echo_tl_state_source,
  input  [1:0]   auto_out_r_bits_echo_extra_id,
  input          auto_out_r_bits_last
);
  assign auto_in_aw_ready = auto_out_aw_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_w_ready = auto_out_w_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_b_valid = auto_out_b_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_b_bits_id = {auto_out_b_bits_echo_extra_id,auto_out_b_bits_id}; // @[Cat.scala 33:92]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_b_bits_echo_tl_state_source = auto_out_b_bits_echo_tl_state_source; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_ar_ready = auto_out_ar_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_valid = auto_out_r_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_bits_id = {auto_out_r_bits_echo_extra_id,auto_out_r_bits_id}; // @[Cat.scala 33:92]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_bits_echo_tl_state_source = auto_out_r_bits_echo_tl_state_source; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_bits_last = auto_out_r_bits_last; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_out_aw_valid = auto_in_aw_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id[5:0]; // @[Nodes.scala 1212:84 BundleMap.scala 247:19]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_len = auto_in_aw_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_size = auto_in_aw_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_burst = auto_in_aw_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_lock = auto_in_aw_bits_lock; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_cache = auto_in_aw_bits_cache; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_prot = auto_in_aw_bits_prot; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_qos = auto_in_aw_bits_qos; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_echo_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_echo_extra_id = auto_in_aw_bits_id[7:6]; // @[IdIndexer.scala 74:56]
  assign auto_out_w_valid = auto_in_w_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_w_bits_strb = auto_in_w_bits_strb; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_b_ready = auto_in_b_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_valid = auto_in_ar_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id[5:0]; // @[Nodes.scala 1212:84 BundleMap.scala 247:19]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_len = auto_in_ar_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_burst = auto_in_ar_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_lock = auto_in_ar_bits_lock; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_cache = auto_in_ar_bits_cache; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_prot = auto_in_ar_bits_prot; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_qos = auto_in_ar_bits_qos; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_echo_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_echo_extra_id = auto_in_ar_bits_id[7:6]; // @[IdIndexer.scala 73:56]
  assign auto_out_r_ready = auto_in_r_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
endmodule
module Queue_166(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [7:0]  io_enq_bits_id,
  input  [33:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_len,
  input  [2:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_burst,
  input         io_enq_bits_lock,
  input  [3:0]  io_enq_bits_cache,
  input  [2:0]  io_enq_bits_prot,
  input  [3:0]  io_enq_bits_qos,
  input  [6:0]  io_enq_bits_echo_tl_state_source,
  input         io_deq_ready,
  output        io_deq_valid,
  output [7:0]  io_deq_bits_id,
  output [33:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_len,
  output [2:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_burst,
  output        io_deq_bits_lock,
  output [3:0]  io_deq_bits_cache,
  output [2:0]  io_deq_bits_prot,
  output [3:0]  io_deq_bits_qos,
  output [6:0]  io_deq_bits_echo_tl_state_source
);
  reg [7:0] ram_id [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [7:0] ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [7:0] ram_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [33:0] ram_addr [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_addr_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_addr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [33:0] ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [33:0] ram_addr_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_addr_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_addr_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_addr_MPORT_en; // @[Decoupled.scala 273:95]
  reg [7:0] ram_len [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_len_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_len_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [7:0] ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [7:0] ram_len_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_len_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_len_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_len_MPORT_en; // @[Decoupled.scala 273:95]
  reg [2:0] ram_size [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_size_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_burst [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_burst_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_burst_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_burst_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_burst_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_burst_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_burst_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_lock [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_lock_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_lock_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_lock_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_lock_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_lock_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_lock_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_lock_MPORT_en; // @[Decoupled.scala 273:95]
  reg [3:0] ram_cache [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_cache_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_cache_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [3:0] ram_cache_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [3:0] ram_cache_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_cache_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_cache_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_cache_MPORT_en; // @[Decoupled.scala 273:95]
  reg [2:0] ram_prot [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_prot_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_prot_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [2:0] ram_prot_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_prot_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_prot_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_prot_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_prot_MPORT_en; // @[Decoupled.scala 273:95]
  reg [3:0] ram_qos [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_qos_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_qos_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [3:0] ram_qos_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [3:0] ram_qos_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_qos_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_qos_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_qos_MPORT_en; // @[Decoupled.scala 273:95]
  reg [6:0] ram_echo_tl_state_source [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [6:0] ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [6:0] ram_echo_tl_state_source_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = enq_ptr_value;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_addr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_addr_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = enq_ptr_value;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_len_io_deq_bits_MPORT_en = 1'h1;
  assign ram_len_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_len_io_deq_bits_MPORT_data = ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_len_MPORT_data = io_enq_bits_len;
  assign ram_len_MPORT_addr = enq_ptr_value;
  assign ram_len_MPORT_mask = 1'h1;
  assign ram_len_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = enq_ptr_value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_burst_io_deq_bits_MPORT_en = 1'h1;
  assign ram_burst_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_burst_io_deq_bits_MPORT_data = ram_burst[ram_burst_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_burst_MPORT_data = io_enq_bits_burst;
  assign ram_burst_MPORT_addr = enq_ptr_value;
  assign ram_burst_MPORT_mask = 1'h1;
  assign ram_burst_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_lock_io_deq_bits_MPORT_en = 1'h1;
  assign ram_lock_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_lock_io_deq_bits_MPORT_data = ram_lock[ram_lock_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_lock_MPORT_data = io_enq_bits_lock;
  assign ram_lock_MPORT_addr = enq_ptr_value;
  assign ram_lock_MPORT_mask = 1'h1;
  assign ram_lock_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_cache_io_deq_bits_MPORT_en = 1'h1;
  assign ram_cache_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_cache_io_deq_bits_MPORT_data = ram_cache[ram_cache_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_cache_MPORT_data = io_enq_bits_cache;
  assign ram_cache_MPORT_addr = enq_ptr_value;
  assign ram_cache_MPORT_mask = 1'h1;
  assign ram_cache_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_prot_io_deq_bits_MPORT_en = 1'h1;
  assign ram_prot_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_prot_io_deq_bits_MPORT_data = ram_prot[ram_prot_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_prot_MPORT_data = io_enq_bits_prot;
  assign ram_prot_MPORT_addr = enq_ptr_value;
  assign ram_prot_MPORT_mask = 1'h1;
  assign ram_prot_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_qos_io_deq_bits_MPORT_en = 1'h1;
  assign ram_qos_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_qos_io_deq_bits_MPORT_data = ram_qos[ram_qos_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_qos_MPORT_data = io_enq_bits_qos;
  assign ram_qos_MPORT_addr = enq_ptr_value;
  assign ram_qos_MPORT_mask = 1'h1;
  assign ram_qos_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_data =
    ram_echo_tl_state_source[ram_echo_tl_state_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_echo_tl_state_source_MPORT_data = io_enq_bits_echo_tl_state_source;
  assign ram_echo_tl_state_source_MPORT_addr = enq_ptr_value;
  assign ram_echo_tl_state_source_MPORT_mask = 1'h1;
  assign ram_echo_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_id = ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_addr = ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_len = ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_burst = ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_lock = ram_lock_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_cache = ram_cache_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_prot = ram_prot_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_qos = ram_qos_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_echo_tl_state_source = ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_len_MPORT_en & ram_len_MPORT_mask) begin
      ram_len[ram_len_MPORT_addr] <= ram_len_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_burst_MPORT_en & ram_burst_MPORT_mask) begin
      ram_burst[ram_burst_MPORT_addr] <= ram_burst_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_lock_MPORT_en & ram_lock_MPORT_mask) begin
      ram_lock[ram_lock_MPORT_addr] <= ram_lock_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_cache_MPORT_en & ram_cache_MPORT_mask) begin
      ram_cache[ram_cache_MPORT_addr] <= ram_cache_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_prot_MPORT_en & ram_prot_MPORT_mask) begin
      ram_prot[ram_prot_MPORT_addr] <= ram_prot_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_qos_MPORT_en & ram_qos_MPORT_mask) begin
      ram_qos[ram_qos_MPORT_addr] <= ram_qos_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_echo_tl_state_source_MPORT_en & ram_echo_tl_state_source_MPORT_mask) begin
      ram_echo_tl_state_source[ram_echo_tl_state_source_MPORT_addr] <= ram_echo_tl_state_source_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
endmodule
module Queue_168(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits_id,
  input  [1:0] io_enq_bits_resp,
  input  [6:0] io_enq_bits_echo_tl_state_source,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits_id,
  output [1:0] io_deq_bits_resp,
  output [6:0] io_deq_bits_echo_tl_state_source
);
  reg [7:0] ram_id [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [7:0] ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [7:0] ram_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_resp [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_resp_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_resp_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_resp_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_en; // @[Decoupled.scala 273:95]
  reg [6:0] ram_echo_tl_state_source [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [6:0] ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [6:0] ram_echo_tl_state_source_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = enq_ptr_value;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_resp_io_deq_bits_MPORT_en = 1'h1;
  assign ram_resp_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_resp_io_deq_bits_MPORT_data = ram_resp[ram_resp_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_resp_MPORT_data = io_enq_bits_resp;
  assign ram_resp_MPORT_addr = enq_ptr_value;
  assign ram_resp_MPORT_mask = 1'h1;
  assign ram_resp_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_data =
    ram_echo_tl_state_source[ram_echo_tl_state_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_echo_tl_state_source_MPORT_data = io_enq_bits_echo_tl_state_source;
  assign ram_echo_tl_state_source_MPORT_addr = enq_ptr_value;
  assign ram_echo_tl_state_source_MPORT_mask = 1'h1;
  assign ram_echo_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_id = ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_resp = ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_echo_tl_state_source = ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_resp_MPORT_en & ram_resp_MPORT_mask) begin
      ram_resp[ram_resp_MPORT_addr] <= ram_resp_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_echo_tl_state_source_MPORT_en & ram_echo_tl_state_source_MPORT_mask) begin
      ram_echo_tl_state_source[ram_echo_tl_state_source_MPORT_addr] <= ram_echo_tl_state_source_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
endmodule
module Queue_170(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [7:0]   io_enq_bits_id,
  input  [511:0] io_enq_bits_data,
  input  [1:0]   io_enq_bits_resp,
  input  [6:0]   io_enq_bits_echo_tl_state_source,
  input          io_enq_bits_last,
  input          io_deq_ready,
  output         io_deq_valid,
  output [7:0]   io_deq_bits_id,
  output [511:0] io_deq_bits_data,
  output [1:0]   io_deq_bits_resp,
  output [6:0]   io_deq_bits_echo_tl_state_source,
  output         io_deq_bits_last
);
  reg [7:0] ram_id [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [7:0] ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [7:0] ram_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [511:0] ram_data [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [511:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [511:0] ram_data_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_resp [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_resp_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_resp_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_resp_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_en; // @[Decoupled.scala 273:95]
  reg [6:0] ram_echo_tl_state_source [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [6:0] ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [6:0] ram_echo_tl_state_source_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_echo_tl_state_source_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_last [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = enq_ptr_value;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_resp_io_deq_bits_MPORT_en = 1'h1;
  assign ram_resp_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_resp_io_deq_bits_MPORT_data = ram_resp[ram_resp_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_resp_MPORT_data = io_enq_bits_resp;
  assign ram_resp_MPORT_addr = enq_ptr_value;
  assign ram_resp_MPORT_mask = 1'h1;
  assign ram_resp_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_data =
    ram_echo_tl_state_source[ram_echo_tl_state_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_echo_tl_state_source_MPORT_data = io_enq_bits_echo_tl_state_source;
  assign ram_echo_tl_state_source_MPORT_addr = enq_ptr_value;
  assign ram_echo_tl_state_source_MPORT_mask = 1'h1;
  assign ram_echo_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_last_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_last_io_deq_bits_MPORT_data = ram_last[ram_last_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_last_MPORT_data = io_enq_bits_last;
  assign ram_last_MPORT_addr = enq_ptr_value;
  assign ram_last_MPORT_mask = 1'h1;
  assign ram_last_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_id = ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_resp = ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_echo_tl_state_source = ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_last = ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_resp_MPORT_en & ram_resp_MPORT_mask) begin
      ram_resp[ram_resp_MPORT_addr] <= ram_resp_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_echo_tl_state_source_MPORT_en & ram_echo_tl_state_source_MPORT_mask) begin
      ram_echo_tl_state_source[ram_echo_tl_state_source_MPORT_addr] <= ram_echo_tl_state_source_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_last_MPORT_en & ram_last_MPORT_mask) begin
      ram_last[ram_last_MPORT_addr] <= ram_last_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
endmodule
module AXI4Buffer_5(
  input          clock,
  input          reset,
  output         auto_in_aw_ready,
  input          auto_in_aw_valid,
  input  [7:0]   auto_in_aw_bits_id,
  input  [33:0]  auto_in_aw_bits_addr,
  input  [7:0]   auto_in_aw_bits_len,
  input  [2:0]   auto_in_aw_bits_size,
  input  [1:0]   auto_in_aw_bits_burst,
  input          auto_in_aw_bits_lock,
  input  [3:0]   auto_in_aw_bits_cache,
  input  [2:0]   auto_in_aw_bits_prot,
  input  [3:0]   auto_in_aw_bits_qos,
  input  [6:0]   auto_in_aw_bits_echo_tl_state_source,
  output         auto_in_w_ready,
  input          auto_in_w_valid,
  input  [511:0] auto_in_w_bits_data,
  input  [63:0]  auto_in_w_bits_strb,
  input          auto_in_w_bits_last,
  input          auto_in_b_ready,
  output         auto_in_b_valid,
  output [7:0]   auto_in_b_bits_id,
  output [1:0]   auto_in_b_bits_resp,
  output [6:0]   auto_in_b_bits_echo_tl_state_source,
  output         auto_in_ar_ready,
  input          auto_in_ar_valid,
  input  [7:0]   auto_in_ar_bits_id,
  input  [33:0]  auto_in_ar_bits_addr,
  input  [7:0]   auto_in_ar_bits_len,
  input  [2:0]   auto_in_ar_bits_size,
  input  [1:0]   auto_in_ar_bits_burst,
  input          auto_in_ar_bits_lock,
  input  [3:0]   auto_in_ar_bits_cache,
  input  [2:0]   auto_in_ar_bits_prot,
  input  [3:0]   auto_in_ar_bits_qos,
  input  [6:0]   auto_in_ar_bits_echo_tl_state_source,
  input          auto_in_r_ready,
  output         auto_in_r_valid,
  output [7:0]   auto_in_r_bits_id,
  output [511:0] auto_in_r_bits_data,
  output [1:0]   auto_in_r_bits_resp,
  output [6:0]   auto_in_r_bits_echo_tl_state_source,
  output         auto_in_r_bits_last,
  input          auto_out_aw_ready,
  output         auto_out_aw_valid,
  output [7:0]   auto_out_aw_bits_id,
  output [33:0]  auto_out_aw_bits_addr,
  output [7:0]   auto_out_aw_bits_len,
  output [2:0]   auto_out_aw_bits_size,
  output [1:0]   auto_out_aw_bits_burst,
  output         auto_out_aw_bits_lock,
  output [3:0]   auto_out_aw_bits_cache,
  output [2:0]   auto_out_aw_bits_prot,
  output [3:0]   auto_out_aw_bits_qos,
  output [6:0]   auto_out_aw_bits_echo_tl_state_source,
  input          auto_out_w_ready,
  output         auto_out_w_valid,
  output [511:0] auto_out_w_bits_data,
  output [63:0]  auto_out_w_bits_strb,
  output         auto_out_w_bits_last,
  output         auto_out_b_ready,
  input          auto_out_b_valid,
  input  [7:0]   auto_out_b_bits_id,
  input  [1:0]   auto_out_b_bits_resp,
  input  [6:0]   auto_out_b_bits_echo_tl_state_source,
  input          auto_out_ar_ready,
  output         auto_out_ar_valid,
  output [7:0]   auto_out_ar_bits_id,
  output [33:0]  auto_out_ar_bits_addr,
  output [7:0]   auto_out_ar_bits_len,
  output [2:0]   auto_out_ar_bits_size,
  output [1:0]   auto_out_ar_bits_burst,
  output         auto_out_ar_bits_lock,
  output [3:0]   auto_out_ar_bits_cache,
  output [2:0]   auto_out_ar_bits_prot,
  output [3:0]   auto_out_ar_bits_qos,
  output [6:0]   auto_out_ar_bits_echo_tl_state_source,
  output         auto_out_r_ready,
  input          auto_out_r_valid,
  input  [7:0]   auto_out_r_bits_id,
  input  [511:0] auto_out_r_bits_data,
  input  [1:0]   auto_out_r_bits_resp,
  input  [6:0]   auto_out_r_bits_echo_tl_state_source,
  input          auto_out_r_bits_last
);
  wire  x1_aw_deq_clock; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_reset; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [7:0] x1_aw_deq_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire [33:0] x1_aw_deq_io_enq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] x1_aw_deq_io_enq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] x1_aw_deq_io_enq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] x1_aw_deq_io_enq_bits_burst; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_enq_bits_lock; // @[Decoupled.scala 375:21]
  wire [3:0] x1_aw_deq_io_enq_bits_cache; // @[Decoupled.scala 375:21]
  wire [2:0] x1_aw_deq_io_enq_bits_prot; // @[Decoupled.scala 375:21]
  wire [3:0] x1_aw_deq_io_enq_bits_qos; // @[Decoupled.scala 375:21]
  wire [6:0] x1_aw_deq_io_enq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [7:0] x1_aw_deq_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [33:0] x1_aw_deq_io_deq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] x1_aw_deq_io_deq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] x1_aw_deq_io_deq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] x1_aw_deq_io_deq_bits_burst; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_deq_bits_lock; // @[Decoupled.scala 375:21]
  wire [3:0] x1_aw_deq_io_deq_bits_cache; // @[Decoupled.scala 375:21]
  wire [2:0] x1_aw_deq_io_deq_bits_prot; // @[Decoupled.scala 375:21]
  wire [3:0] x1_aw_deq_io_deq_bits_qos; // @[Decoupled.scala 375:21]
  wire [6:0] x1_aw_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_clock; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_reset; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [511:0] x1_w_deq_io_enq_bits_data; // @[Decoupled.scala 375:21]
  wire [63:0] x1_w_deq_io_enq_bits_strb; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_enq_bits_last; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [511:0] x1_w_deq_io_deq_bits_data; // @[Decoupled.scala 375:21]
  wire [63:0] x1_w_deq_io_deq_bits_strb; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_deq_bits_last; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_clock; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_reset; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [7:0] bundleIn_0_b_deq_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire [1:0] bundleIn_0_b_deq_io_enq_bits_resp; // @[Decoupled.scala 375:21]
  wire [6:0] bundleIn_0_b_deq_io_enq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [7:0] bundleIn_0_b_deq_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [1:0] bundleIn_0_b_deq_io_deq_bits_resp; // @[Decoupled.scala 375:21]
  wire [6:0] bundleIn_0_b_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_clock; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_reset; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [7:0] x1_ar_deq_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire [33:0] x1_ar_deq_io_enq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] x1_ar_deq_io_enq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] x1_ar_deq_io_enq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] x1_ar_deq_io_enq_bits_burst; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_enq_bits_lock; // @[Decoupled.scala 375:21]
  wire [3:0] x1_ar_deq_io_enq_bits_cache; // @[Decoupled.scala 375:21]
  wire [2:0] x1_ar_deq_io_enq_bits_prot; // @[Decoupled.scala 375:21]
  wire [3:0] x1_ar_deq_io_enq_bits_qos; // @[Decoupled.scala 375:21]
  wire [6:0] x1_ar_deq_io_enq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [7:0] x1_ar_deq_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [33:0] x1_ar_deq_io_deq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] x1_ar_deq_io_deq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] x1_ar_deq_io_deq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] x1_ar_deq_io_deq_bits_burst; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_deq_bits_lock; // @[Decoupled.scala 375:21]
  wire [3:0] x1_ar_deq_io_deq_bits_cache; // @[Decoupled.scala 375:21]
  wire [2:0] x1_ar_deq_io_deq_bits_prot; // @[Decoupled.scala 375:21]
  wire [3:0] x1_ar_deq_io_deq_bits_qos; // @[Decoupled.scala 375:21]
  wire [6:0] x1_ar_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_clock; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_reset; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [7:0] bundleIn_0_r_deq_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire [511:0] bundleIn_0_r_deq_io_enq_bits_data; // @[Decoupled.scala 375:21]
  wire [1:0] bundleIn_0_r_deq_io_enq_bits_resp; // @[Decoupled.scala 375:21]
  wire [6:0] bundleIn_0_r_deq_io_enq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_enq_bits_last; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [7:0] bundleIn_0_r_deq_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [511:0] bundleIn_0_r_deq_io_deq_bits_data; // @[Decoupled.scala 375:21]
  wire [1:0] bundleIn_0_r_deq_io_deq_bits_resp; // @[Decoupled.scala 375:21]
  wire [6:0] bundleIn_0_r_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_deq_bits_last; // @[Decoupled.scala 375:21]
  Queue_166 x1_aw_deq ( // @[Decoupled.scala 375:21]
    .clock(x1_aw_deq_clock),
    .reset(x1_aw_deq_reset),
    .io_enq_ready(x1_aw_deq_io_enq_ready),
    .io_enq_valid(x1_aw_deq_io_enq_valid),
    .io_enq_bits_id(x1_aw_deq_io_enq_bits_id),
    .io_enq_bits_addr(x1_aw_deq_io_enq_bits_addr),
    .io_enq_bits_len(x1_aw_deq_io_enq_bits_len),
    .io_enq_bits_size(x1_aw_deq_io_enq_bits_size),
    .io_enq_bits_burst(x1_aw_deq_io_enq_bits_burst),
    .io_enq_bits_lock(x1_aw_deq_io_enq_bits_lock),
    .io_enq_bits_cache(x1_aw_deq_io_enq_bits_cache),
    .io_enq_bits_prot(x1_aw_deq_io_enq_bits_prot),
    .io_enq_bits_qos(x1_aw_deq_io_enq_bits_qos),
    .io_enq_bits_echo_tl_state_source(x1_aw_deq_io_enq_bits_echo_tl_state_source),
    .io_deq_ready(x1_aw_deq_io_deq_ready),
    .io_deq_valid(x1_aw_deq_io_deq_valid),
    .io_deq_bits_id(x1_aw_deq_io_deq_bits_id),
    .io_deq_bits_addr(x1_aw_deq_io_deq_bits_addr),
    .io_deq_bits_len(x1_aw_deq_io_deq_bits_len),
    .io_deq_bits_size(x1_aw_deq_io_deq_bits_size),
    .io_deq_bits_burst(x1_aw_deq_io_deq_bits_burst),
    .io_deq_bits_lock(x1_aw_deq_io_deq_bits_lock),
    .io_deq_bits_cache(x1_aw_deq_io_deq_bits_cache),
    .io_deq_bits_prot(x1_aw_deq_io_deq_bits_prot),
    .io_deq_bits_qos(x1_aw_deq_io_deq_bits_qos),
    .io_deq_bits_echo_tl_state_source(x1_aw_deq_io_deq_bits_echo_tl_state_source)
  );
  Queue_7 x1_w_deq ( // @[Decoupled.scala 375:21]
    .clock(x1_w_deq_clock),
    .reset(x1_w_deq_reset),
    .io_enq_ready(x1_w_deq_io_enq_ready),
    .io_enq_valid(x1_w_deq_io_enq_valid),
    .io_enq_bits_data(x1_w_deq_io_enq_bits_data),
    .io_enq_bits_strb(x1_w_deq_io_enq_bits_strb),
    .io_enq_bits_last(x1_w_deq_io_enq_bits_last),
    .io_deq_ready(x1_w_deq_io_deq_ready),
    .io_deq_valid(x1_w_deq_io_deq_valid),
    .io_deq_bits_data(x1_w_deq_io_deq_bits_data),
    .io_deq_bits_strb(x1_w_deq_io_deq_bits_strb),
    .io_deq_bits_last(x1_w_deq_io_deq_bits_last)
  );
  Queue_168 bundleIn_0_b_deq ( // @[Decoupled.scala 375:21]
    .clock(bundleIn_0_b_deq_clock),
    .reset(bundleIn_0_b_deq_reset),
    .io_enq_ready(bundleIn_0_b_deq_io_enq_ready),
    .io_enq_valid(bundleIn_0_b_deq_io_enq_valid),
    .io_enq_bits_id(bundleIn_0_b_deq_io_enq_bits_id),
    .io_enq_bits_resp(bundleIn_0_b_deq_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_source(bundleIn_0_b_deq_io_enq_bits_echo_tl_state_source),
    .io_deq_ready(bundleIn_0_b_deq_io_deq_ready),
    .io_deq_valid(bundleIn_0_b_deq_io_deq_valid),
    .io_deq_bits_id(bundleIn_0_b_deq_io_deq_bits_id),
    .io_deq_bits_resp(bundleIn_0_b_deq_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_source(bundleIn_0_b_deq_io_deq_bits_echo_tl_state_source)
  );
  Queue_166 x1_ar_deq ( // @[Decoupled.scala 375:21]
    .clock(x1_ar_deq_clock),
    .reset(x1_ar_deq_reset),
    .io_enq_ready(x1_ar_deq_io_enq_ready),
    .io_enq_valid(x1_ar_deq_io_enq_valid),
    .io_enq_bits_id(x1_ar_deq_io_enq_bits_id),
    .io_enq_bits_addr(x1_ar_deq_io_enq_bits_addr),
    .io_enq_bits_len(x1_ar_deq_io_enq_bits_len),
    .io_enq_bits_size(x1_ar_deq_io_enq_bits_size),
    .io_enq_bits_burst(x1_ar_deq_io_enq_bits_burst),
    .io_enq_bits_lock(x1_ar_deq_io_enq_bits_lock),
    .io_enq_bits_cache(x1_ar_deq_io_enq_bits_cache),
    .io_enq_bits_prot(x1_ar_deq_io_enq_bits_prot),
    .io_enq_bits_qos(x1_ar_deq_io_enq_bits_qos),
    .io_enq_bits_echo_tl_state_source(x1_ar_deq_io_enq_bits_echo_tl_state_source),
    .io_deq_ready(x1_ar_deq_io_deq_ready),
    .io_deq_valid(x1_ar_deq_io_deq_valid),
    .io_deq_bits_id(x1_ar_deq_io_deq_bits_id),
    .io_deq_bits_addr(x1_ar_deq_io_deq_bits_addr),
    .io_deq_bits_len(x1_ar_deq_io_deq_bits_len),
    .io_deq_bits_size(x1_ar_deq_io_deq_bits_size),
    .io_deq_bits_burst(x1_ar_deq_io_deq_bits_burst),
    .io_deq_bits_lock(x1_ar_deq_io_deq_bits_lock),
    .io_deq_bits_cache(x1_ar_deq_io_deq_bits_cache),
    .io_deq_bits_prot(x1_ar_deq_io_deq_bits_prot),
    .io_deq_bits_qos(x1_ar_deq_io_deq_bits_qos),
    .io_deq_bits_echo_tl_state_source(x1_ar_deq_io_deq_bits_echo_tl_state_source)
  );
  Queue_170 bundleIn_0_r_deq ( // @[Decoupled.scala 375:21]
    .clock(bundleIn_0_r_deq_clock),
    .reset(bundleIn_0_r_deq_reset),
    .io_enq_ready(bundleIn_0_r_deq_io_enq_ready),
    .io_enq_valid(bundleIn_0_r_deq_io_enq_valid),
    .io_enq_bits_id(bundleIn_0_r_deq_io_enq_bits_id),
    .io_enq_bits_data(bundleIn_0_r_deq_io_enq_bits_data),
    .io_enq_bits_resp(bundleIn_0_r_deq_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_source(bundleIn_0_r_deq_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(bundleIn_0_r_deq_io_enq_bits_last),
    .io_deq_ready(bundleIn_0_r_deq_io_deq_ready),
    .io_deq_valid(bundleIn_0_r_deq_io_deq_valid),
    .io_deq_bits_id(bundleIn_0_r_deq_io_deq_bits_id),
    .io_deq_bits_data(bundleIn_0_r_deq_io_deq_bits_data),
    .io_deq_bits_resp(bundleIn_0_r_deq_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_source(bundleIn_0_r_deq_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(bundleIn_0_r_deq_io_deq_bits_last)
  );
  assign auto_in_aw_ready = x1_aw_deq_io_enq_ready; // @[Nodes.scala 1215:84 Decoupled.scala 379:17]
  assign auto_in_w_ready = x1_w_deq_io_enq_ready; // @[Nodes.scala 1215:84 Decoupled.scala 379:17]
  assign auto_in_b_valid = bundleIn_0_b_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_in_b_bits_id = bundleIn_0_b_deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_b_bits_resp = bundleIn_0_b_deq_io_deq_bits_resp; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_b_bits_echo_tl_state_source = bundleIn_0_b_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_ar_ready = x1_ar_deq_io_enq_ready; // @[Nodes.scala 1215:84 Decoupled.scala 379:17]
  assign auto_in_r_valid = bundleIn_0_r_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_in_r_bits_id = bundleIn_0_r_deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_r_bits_data = bundleIn_0_r_deq_io_deq_bits_data; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_r_bits_resp = bundleIn_0_r_deq_io_deq_bits_resp; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_r_bits_echo_tl_state_source = bundleIn_0_r_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_r_bits_last = bundleIn_0_r_deq_io_deq_bits_last; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_valid = x1_aw_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_out_aw_bits_id = x1_aw_deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_addr = x1_aw_deq_io_deq_bits_addr; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_len = x1_aw_deq_io_deq_bits_len; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_size = x1_aw_deq_io_deq_bits_size; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_burst = x1_aw_deq_io_deq_bits_burst; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_lock = x1_aw_deq_io_deq_bits_lock; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_cache = x1_aw_deq_io_deq_bits_cache; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_prot = x1_aw_deq_io_deq_bits_prot; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_qos = x1_aw_deq_io_deq_bits_qos; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_echo_tl_state_source = x1_aw_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_w_valid = x1_w_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_out_w_bits_data = x1_w_deq_io_deq_bits_data; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_w_bits_strb = x1_w_deq_io_deq_bits_strb; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_w_bits_last = x1_w_deq_io_deq_bits_last; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_b_ready = bundleIn_0_b_deq_io_enq_ready; // @[Nodes.scala 1212:84 Decoupled.scala 379:17]
  assign auto_out_ar_valid = x1_ar_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_out_ar_bits_id = x1_ar_deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_addr = x1_ar_deq_io_deq_bits_addr; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_len = x1_ar_deq_io_deq_bits_len; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_size = x1_ar_deq_io_deq_bits_size; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_burst = x1_ar_deq_io_deq_bits_burst; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_lock = x1_ar_deq_io_deq_bits_lock; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_cache = x1_ar_deq_io_deq_bits_cache; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_prot = x1_ar_deq_io_deq_bits_prot; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_qos = x1_ar_deq_io_deq_bits_qos; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_echo_tl_state_source = x1_ar_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_r_ready = bundleIn_0_r_deq_io_enq_ready; // @[Nodes.scala 1212:84 Decoupled.scala 379:17]
  assign x1_aw_deq_clock = clock;
  assign x1_aw_deq_reset = reset;
  assign x1_aw_deq_io_enq_valid = auto_in_aw_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_id = auto_in_aw_bits_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_addr = auto_in_aw_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_len = auto_in_aw_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_size = auto_in_aw_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_burst = auto_in_aw_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_lock = auto_in_aw_bits_lock; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_cache = auto_in_aw_bits_cache; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_prot = auto_in_aw_bits_prot; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_qos = auto_in_aw_bits_qos; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_echo_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_deq_ready = auto_out_aw_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign x1_w_deq_clock = clock;
  assign x1_w_deq_reset = reset;
  assign x1_w_deq_io_enq_valid = auto_in_w_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_w_deq_io_enq_bits_data = auto_in_w_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_w_deq_io_enq_bits_strb = auto_in_w_bits_strb; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_w_deq_io_enq_bits_last = auto_in_w_bits_last; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_w_deq_io_deq_ready = auto_out_w_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_b_deq_clock = clock;
  assign bundleIn_0_b_deq_reset = reset;
  assign bundleIn_0_b_deq_io_enq_valid = auto_out_b_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_b_deq_io_enq_bits_id = auto_out_b_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_b_deq_io_enq_bits_resp = auto_out_b_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_b_deq_io_enq_bits_echo_tl_state_source = auto_out_b_bits_echo_tl_state_source; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_b_deq_io_deq_ready = auto_in_b_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_clock = clock;
  assign x1_ar_deq_reset = reset;
  assign x1_ar_deq_io_enq_valid = auto_in_ar_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_id = auto_in_ar_bits_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_addr = auto_in_ar_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_len = auto_in_ar_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_size = auto_in_ar_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_burst = auto_in_ar_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_lock = auto_in_ar_bits_lock; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_cache = auto_in_ar_bits_cache; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_prot = auto_in_ar_bits_prot; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_qos = auto_in_ar_bits_qos; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_echo_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_deq_ready = auto_out_ar_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_clock = clock;
  assign bundleIn_0_r_deq_reset = reset;
  assign bundleIn_0_r_deq_io_enq_valid = auto_out_r_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_enq_bits_id = auto_out_r_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_enq_bits_data = auto_out_r_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_enq_bits_resp = auto_out_r_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_enq_bits_echo_tl_state_source = auto_out_r_bits_echo_tl_state_source; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_enq_bits_last = auto_out_r_bits_last; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_deq_ready = auto_in_r_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
endmodule
module MCRFileTL(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [3:0]  auto_in_a_bits_source,
  input  [15:0] auto_in_a_bits_address,
  input  [31:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [3:0]  auto_in_d_bits_source,
  output [31:0] auto_in_d_bits_data,
  output        io_mcr_read_0_ready,
  input  [31:0] io_mcr_read_0_bits,
  output        io_mcr_read_1_ready,
  input  [31:0] io_mcr_read_1_bits,
  output        io_mcr_read_2_ready,
  input  [31:0] io_mcr_read_2_bits,
  output        io_mcr_read_3_ready,
  input  [31:0] io_mcr_read_3_bits,
  output        io_mcr_read_4_ready,
  input  [31:0] io_mcr_read_4_bits,
  output        io_mcr_read_5_ready,
  input  [31:0] io_mcr_read_5_bits,
  output        io_mcr_read_6_ready,
  input  [31:0] io_mcr_read_6_bits,
  output        io_mcr_read_7_ready,
  output        io_mcr_write_0_valid,
  output [31:0] io_mcr_write_0_bits,
  output        io_mcr_write_1_valid,
  output [31:0] io_mcr_write_1_bits,
  output        io_mcr_write_2_valid,
  output [31:0] io_mcr_write_2_bits,
  output        io_mcr_write_3_valid,
  output [31:0] io_mcr_write_3_bits,
  output        io_mcr_write_4_valid,
  output [31:0] io_mcr_write_4_bits,
  output        io_mcr_write_5_valid,
  output [31:0] io_mcr_write_5_bits,
  output        io_mcr_write_6_valid,
  output [31:0] io_mcr_write_6_bits
);
  reg [2:0] state; // @[MCR.scala 268:22]
  reg [2:0] address; // @[MCR.scala 270:20]
  reg [31:0] writeData; // @[MCR.scala 271:22]
  reg [31:0] readData; // @[MCR.scala 272:21]
  reg [3:0] id; // @[MCR.scala 273:15]
  wire  in_a_ready = 3'h0 == state; // @[MCR.scala 292:17]
  wire  _T_1 = in_a_ready & auto_in_a_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_0 = auto_in_a_bits_opcode == 3'h0 | auto_in_a_bits_opcode == 3'h1 ? 3'h3 : state; // @[MCR.scala 302:110 303:17 268:22]
  wire  _GEN_16 = 3'h0 == address; // @[MCR.scala 284:20 313:{35,35}]
  wire  _GEN_17 = 3'h1 == address; // @[MCR.scala 284:20 313:{35,35}]
  wire  _GEN_18 = 3'h2 == address; // @[MCR.scala 284:20 313:{35,35}]
  wire  _GEN_19 = 3'h3 == address; // @[MCR.scala 284:20 313:{35,35}]
  wire  _GEN_20 = 3'h4 == address; // @[MCR.scala 284:20 313:{35,35}]
  wire  _GEN_21 = 3'h5 == address; // @[MCR.scala 284:20 313:{35,35}]
  wire  _GEN_22 = 3'h6 == address; // @[MCR.scala 284:20 313:{35,35}]
  wire  _GEN_23 = 3'h7 == address; // @[MCR.scala 284:20 313:{35,35}]
  wire  _GEN_79 = 3'h1 == state ? 1'h0 : 3'h2 == state; // @[MCR.scala 288:14 292:17]
  wire  _GEN_88 = 3'h4 == state | _GEN_79; // @[MCR.scala 292:17 317:18]
  wire  _GEN_124 = 3'h3 == state ? 1'h0 : _GEN_88; // @[MCR.scala 288:14 292:17]
  wire  in_d_valid = in_a_ready ? 1'h0 : _GEN_124; // @[MCR.scala 288:14 292:17]
  wire  _T_8 = auto_in_d_ready & in_d_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_24 = _T_8 ? 3'h0 : state; // @[MCR.scala 319:24 320:15 268:22]
  wire [31:0] _GEN_34 = 3'h1 == address ? io_mcr_read_1_bits : io_mcr_read_0_bits; // @[MCR.scala 325:{16,16}]
  wire [31:0] _GEN_35 = 3'h2 == address ? io_mcr_read_2_bits : _GEN_34; // @[MCR.scala 325:{16,16}]
  wire [31:0] _GEN_36 = 3'h3 == address ? io_mcr_read_3_bits : _GEN_35; // @[MCR.scala 325:{16,16}]
  wire [31:0] _GEN_37 = 3'h4 == address ? io_mcr_read_4_bits : _GEN_36; // @[MCR.scala 325:{16,16}]
  wire [31:0] _GEN_38 = 3'h5 == address ? io_mcr_read_5_bits : _GEN_37; // @[MCR.scala 325:{16,16}]
  wire [31:0] _GEN_39 = 3'h6 == address ? io_mcr_read_6_bits : _GEN_38; // @[MCR.scala 325:{16,16}]
  wire [31:0] _GEN_40 = 3'h7 == address ? 32'h0 : _GEN_39; // @[MCR.scala 325:{16,16}]
  wire  _GEN_42 = 3'h1 == address ? io_mcr_read_1_ready : io_mcr_read_0_ready; // @[Decoupled.scala 51:{35,35}]
  wire  _GEN_43 = 3'h2 == address ? io_mcr_read_2_ready : _GEN_42; // @[Decoupled.scala 51:{35,35}]
  wire  _GEN_44 = 3'h3 == address ? io_mcr_read_3_ready : _GEN_43; // @[Decoupled.scala 51:{35,35}]
  wire  _GEN_45 = 3'h4 == address ? io_mcr_read_4_ready : _GEN_44; // @[Decoupled.scala 51:{35,35}]
  wire  _GEN_46 = 3'h5 == address ? io_mcr_read_5_ready : _GEN_45; // @[Decoupled.scala 51:{35,35}]
  wire  _GEN_47 = 3'h6 == address ? io_mcr_read_6_ready : _GEN_46; // @[Decoupled.scala 51:{35,35}]
  wire  _GEN_48 = 3'h7 == address ? io_mcr_read_7_ready : _GEN_47; // @[Decoupled.scala 51:{35,35}]
  wire  _GEN_56 = 3'h7 == address ? 1'h0 : 1'h1; // @[Decoupled.scala 51:{35,35}]
  wire  _T_10 = _GEN_48 & _GEN_56; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_57 = _T_10 ? 3'h2 : state; // @[MCR.scala 326:39 327:15 268:22]
  wire [2:0] _GEN_68 = 3'h2 == state ? _GEN_24 : state; // @[MCR.scala 292:17 268:22]
  wire [2:0] _GEN_78 = 3'h1 == state ? _GEN_57 : _GEN_68; // @[MCR.scala 292:17]
  wire  _GEN_98 = 3'h4 == state ? 1'h0 : 3'h1 == state & _GEN_16; // @[MCR.scala 292:17 280:20]
  wire  _GEN_99 = 3'h4 == state ? 1'h0 : 3'h1 == state & _GEN_17; // @[MCR.scala 292:17 280:20]
  wire  _GEN_100 = 3'h4 == state ? 1'h0 : 3'h1 == state & _GEN_18; // @[MCR.scala 292:17 280:20]
  wire  _GEN_101 = 3'h4 == state ? 1'h0 : 3'h1 == state & _GEN_19; // @[MCR.scala 292:17 280:20]
  wire  _GEN_102 = 3'h4 == state ? 1'h0 : 3'h1 == state & _GEN_20; // @[MCR.scala 292:17 280:20]
  wire  _GEN_103 = 3'h4 == state ? 1'h0 : 3'h1 == state & _GEN_21; // @[MCR.scala 292:17 280:20]
  wire  _GEN_104 = 3'h4 == state ? 1'h0 : 3'h1 == state & _GEN_22; // @[MCR.scala 292:17 280:20]
  wire  _GEN_105 = 3'h4 == state ? 1'h0 : 3'h1 == state & _GEN_23; // @[MCR.scala 292:17 280:20]
  wire  _GEN_133 = 3'h3 == state ? 1'h0 : _GEN_98; // @[MCR.scala 292:17 280:20]
  wire  _GEN_134 = 3'h3 == state ? 1'h0 : _GEN_99; // @[MCR.scala 292:17 280:20]
  wire  _GEN_135 = 3'h3 == state ? 1'h0 : _GEN_100; // @[MCR.scala 292:17 280:20]
  wire  _GEN_136 = 3'h3 == state ? 1'h0 : _GEN_101; // @[MCR.scala 292:17 280:20]
  wire  _GEN_137 = 3'h3 == state ? 1'h0 : _GEN_102; // @[MCR.scala 292:17 280:20]
  wire  _GEN_138 = 3'h3 == state ? 1'h0 : _GEN_103; // @[MCR.scala 292:17 280:20]
  wire  _GEN_139 = 3'h3 == state ? 1'h0 : _GEN_104; // @[MCR.scala 292:17 280:20]
  wire  _GEN_140 = 3'h3 == state ? 1'h0 : _GEN_105; // @[MCR.scala 292:17 280:20]
  assign auto_in_a_ready = 3'h0 == state; // @[MCR.scala 292:17]
  assign auto_in_d_valid = in_a_ready ? 1'h0 : _GEN_124; // @[MCR.scala 288:14 292:17]
  assign auto_in_d_bits_opcode = 3'h4 == state ? 3'h0 : 3'h1; // @[MCR.scala 292:17 318:17]
  assign auto_in_d_bits_source = id; // @[MCR.scala 292:17 318:17]
  assign auto_in_d_bits_data = 3'h4 == state ? 32'h0 : readData; // @[MCR.scala 292:17 318:17]
  assign io_mcr_read_0_ready = in_a_ready ? 1'h0 : _GEN_133; // @[MCR.scala 292:17 280:20]
  assign io_mcr_read_1_ready = in_a_ready ? 1'h0 : _GEN_134; // @[MCR.scala 292:17 280:20]
  assign io_mcr_read_2_ready = in_a_ready ? 1'h0 : _GEN_135; // @[MCR.scala 292:17 280:20]
  assign io_mcr_read_3_ready = in_a_ready ? 1'h0 : _GEN_136; // @[MCR.scala 292:17 280:20]
  assign io_mcr_read_4_ready = in_a_ready ? 1'h0 : _GEN_137; // @[MCR.scala 292:17 280:20]
  assign io_mcr_read_5_ready = in_a_ready ? 1'h0 : _GEN_138; // @[MCR.scala 292:17 280:20]
  assign io_mcr_read_6_ready = in_a_ready ? 1'h0 : _GEN_139; // @[MCR.scala 292:17 280:20]
  assign io_mcr_read_7_ready = in_a_ready ? 1'h0 : _GEN_140; // @[MCR.scala 292:17 280:20]
  assign io_mcr_write_0_valid = in_a_ready ? 1'h0 : 3'h3 == state & _GEN_16; // @[MCR.scala 292:17 284:20]
  assign io_mcr_write_0_bits = writeData; // @[MCR.scala 312:{34,34}]
  assign io_mcr_write_1_valid = in_a_ready ? 1'h0 : 3'h3 == state & _GEN_17; // @[MCR.scala 292:17 284:20]
  assign io_mcr_write_1_bits = writeData; // @[MCR.scala 312:{34,34}]
  assign io_mcr_write_2_valid = in_a_ready ? 1'h0 : 3'h3 == state & _GEN_18; // @[MCR.scala 292:17 284:20]
  assign io_mcr_write_2_bits = writeData; // @[MCR.scala 312:{34,34}]
  assign io_mcr_write_3_valid = in_a_ready ? 1'h0 : 3'h3 == state & _GEN_19; // @[MCR.scala 292:17 284:20]
  assign io_mcr_write_3_bits = writeData; // @[MCR.scala 312:{34,34}]
  assign io_mcr_write_4_valid = in_a_ready ? 1'h0 : 3'h3 == state & _GEN_20; // @[MCR.scala 292:17 284:20]
  assign io_mcr_write_4_bits = writeData; // @[MCR.scala 312:{34,34}]
  assign io_mcr_write_5_valid = in_a_ready ? 1'h0 : 3'h3 == state & _GEN_21; // @[MCR.scala 292:17 284:20]
  assign io_mcr_write_5_bits = writeData; // @[MCR.scala 312:{34,34}]
  assign io_mcr_write_6_valid = in_a_ready ? 1'h0 : 3'h3 == state & _GEN_22; // @[MCR.scala 292:17 284:20]
  assign io_mcr_write_6_bits = writeData; // @[MCR.scala 312:{34,34}]
  always @(posedge clock) begin
    if (reset) begin // @[MCR.scala 268:22]
      state <= 3'h0; // @[MCR.scala 268:22]
    end else if (in_a_ready) begin // @[MCR.scala 292:17]
      if (_T_1) begin // @[MCR.scala 295:24]
        if (auto_in_a_bits_opcode == 3'h4) begin // @[MCR.scala 306:52]
          state <= 3'h1; // @[MCR.scala 307:17]
        end else begin
          state <= _GEN_0;
        end
      end
    end else if (3'h3 == state) begin // @[MCR.scala 292:17]
      state <= 3'h4; // @[MCR.scala 314:13]
    end else if (3'h4 == state) begin // @[MCR.scala 292:17]
      state <= _GEN_24;
    end else begin
      state <= _GEN_78;
    end
    if (in_a_ready) begin // @[MCR.scala 292:17]
      if (_T_1) begin // @[MCR.scala 295:24]
        address <= auto_in_a_bits_address[4:2]; // @[MCR.scala 301:17]
      end
    end
    if (in_a_ready) begin // @[MCR.scala 292:17]
      if (_T_1) begin // @[MCR.scala 295:24]
        if (auto_in_a_bits_opcode == 3'h0 | auto_in_a_bits_opcode == 3'h1) begin // @[MCR.scala 302:110]
          writeData <= auto_in_a_bits_data; // @[MCR.scala 304:21]
        end
      end
    end
    if (!(in_a_ready)) begin // @[MCR.scala 292:17]
      if (!(3'h3 == state)) begin // @[MCR.scala 292:17]
        if (!(3'h4 == state)) begin // @[MCR.scala 292:17]
          if (3'h1 == state) begin // @[MCR.scala 292:17]
            readData <= _GEN_40; // @[MCR.scala 325:16]
          end
        end
      end
    end
    if (in_a_ready) begin // @[MCR.scala 292:17]
      if (_T_1) begin // @[MCR.scala 295:24]
        id <= auto_in_a_bits_source; // @[MCR.scala 296:12]
      end
    end
  end
endmodule
module Queue_171(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_id,
  input  [31:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_id,
  output [31:0] io_deq_bits_data,
  output [1:0]  io_deq_bits_resp,
  output        io_deq_bits_last
);
  reg  ram_id [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [31:0] ram_data [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [31:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [31:0] ram_data_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_resp [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_resp_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_resp_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_resp_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_last [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_en; // @[Decoupled.scala 273:95]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 278:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_12 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 318:26 280:27 318:35]
  wire  do_enq = empty ? _GEN_12 : _do_enq_T; // @[Decoupled.scala 315:17 280:27]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 315:17 317:14 281:27]
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = 1'h0;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = 1'h0;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign ram_resp_io_deq_bits_MPORT_en = 1'h1;
  assign ram_resp_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_resp_io_deq_bits_MPORT_data = ram_resp[ram_resp_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_resp_MPORT_data = 2'h0;
  assign ram_resp_MPORT_addr = 1'h0;
  assign ram_resp_MPORT_mask = 1'h1;
  assign ram_resp_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign ram_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_last_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_last_io_deq_bits_MPORT_data = ram_last[ram_last_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_last_MPORT_data = 1'h1;
  assign ram_last_MPORT_addr = 1'h0;
  assign ram_last_MPORT_mask = 1'h1;
  assign ram_last_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 302:16 314:{24,39}]
  assign io_deq_bits_id = empty ? io_enq_bits_id : ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_data = empty ? io_enq_bits_data : ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_resp = empty ? 2'h0 : ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_last = empty | ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_resp_MPORT_en & ram_resp_MPORT_mask) begin
      ram_resp[ram_resp_MPORT_addr] <= ram_resp_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_last_MPORT_en & ram_last_MPORT_mask) begin
      ram_last[ram_last_MPORT_addr] <= ram_last_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      if (empty) begin // @[Decoupled.scala 315:17]
        if (io_deq_ready) begin // @[Decoupled.scala 318:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 318:35]
        end else begin
          maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
        end
      end else begin
        maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
      end
    end
  end
endmodule
module Queue_172(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input        io_enq_bits_id,
  input        io_deq_ready,
  output       io_deq_valid,
  output       io_deq_bits_id,
  output [1:0] io_deq_bits_resp
);
  reg  ram_id [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_resp [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_resp_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_resp_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_resp_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_en; // @[Decoupled.scala 273:95]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 278:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_10 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 318:26 280:27 318:35]
  wire  do_enq = empty ? _GEN_10 : _do_enq_T; // @[Decoupled.scala 315:17 280:27]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 315:17 317:14 281:27]
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = 1'h0;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = empty ? _GEN_10 : _do_enq_T;
  assign ram_resp_io_deq_bits_MPORT_en = 1'h1;
  assign ram_resp_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_resp_io_deq_bits_MPORT_data = ram_resp[ram_resp_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_resp_MPORT_data = 2'h0;
  assign ram_resp_MPORT_addr = 1'h0;
  assign ram_resp_MPORT_mask = 1'h1;
  assign ram_resp_MPORT_en = empty ? _GEN_10 : _do_enq_T;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 302:16 314:{24,39}]
  assign io_deq_bits_id = empty ? io_enq_bits_id : ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_resp = empty ? 2'h0 : ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_resp_MPORT_en & ram_resp_MPORT_mask) begin
      ram_resp[ram_resp_MPORT_addr] <= ram_resp_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      if (empty) begin // @[Decoupled.scala 315:17]
        if (io_deq_ready) begin // @[Decoupled.scala 318:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 318:35]
        end else begin
          maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
        end
      end else begin
        maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
      end
    end
  end
endmodule
module AXI4ToTL(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [15:0] auto_in_aw_bits_addr,
  input  [2:0]  auto_in_aw_bits_size,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output        auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [15:0] auto_in_ar_bits_addr,
  input  [2:0]  auto_in_ar_bits_size,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output        auto_in_r_bits_id,
  output [31:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [3:0]  auto_out_a_bits_source,
  output [15:0] auto_out_a_bits_address,
  output [31:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [3:0]  auto_out_d_bits_source,
  input  [31:0] auto_out_d_bits_data
);
  wire  deq_clock; // @[Decoupled.scala 375:21]
  wire  deq_reset; // @[Decoupled.scala 375:21]
  wire  deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire  deq_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire [31:0] deq_io_enq_bits_data; // @[Decoupled.scala 375:21]
  wire  deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire  deq_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [31:0] deq_io_deq_bits_data; // @[Decoupled.scala 375:21]
  wire [1:0] deq_io_deq_bits_resp; // @[Decoupled.scala 375:21]
  wire  deq_io_deq_bits_last; // @[Decoupled.scala 375:21]
  wire  q_b_deq_clock; // @[Decoupled.scala 375:21]
  wire  q_b_deq_reset; // @[Decoupled.scala 375:21]
  wire  q_b_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  q_b_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire  q_b_deq_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire  q_b_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  q_b_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire  q_b_deq_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [1:0] q_b_deq_io_deq_bits_resp; // @[Decoupled.scala 375:21]
  wire [22:0] _r_size1_T_1 = 23'hff << auto_in_ar_bits_size; // @[Bundles.scala 33:21]
  wire [14:0] r_size1 = _r_size1_T_1[22:8]; // @[Bundles.scala 33:30]
  wire [15:0] _r_size_T = {r_size1, 1'h0}; // @[package.scala 233:35]
  wire [15:0] _r_size_T_1 = _r_size_T | 16'h1; // @[package.scala 233:40]
  wire [15:0] _r_size_T_2 = {1'h0,r_size1}; // @[Cat.scala 33:92]
  wire [15:0] _r_size_T_3 = ~_r_size_T_2; // @[package.scala 233:49]
  wire [15:0] _r_size_T_4 = _r_size_T_1 & _r_size_T_3; // @[package.scala 233:47]
  wire [7:0] r_size_hi = _r_size_T_4[15:8]; // @[OneHot.scala 30:18]
  wire [7:0] r_size_lo = _r_size_T_4[7:0]; // @[OneHot.scala 31:18]
  wire  _r_size_T_5 = |r_size_hi; // @[OneHot.scala 32:14]
  wire [7:0] _r_size_T_6 = r_size_hi | r_size_lo; // @[OneHot.scala 32:28]
  wire [3:0] r_size_hi_1 = _r_size_T_6[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] r_size_lo_1 = _r_size_T_6[3:0]; // @[OneHot.scala 31:18]
  wire  _r_size_T_7 = |r_size_hi_1; // @[OneHot.scala 32:14]
  wire [3:0] _r_size_T_8 = r_size_hi_1 | r_size_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] r_size_hi_2 = _r_size_T_8[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] r_size_lo_2 = _r_size_T_8[1:0]; // @[OneHot.scala 31:18]
  wire  _r_size_T_9 = |r_size_hi_2; // @[OneHot.scala 32:14]
  wire [1:0] _r_size_T_10 = r_size_hi_2 | r_size_lo_2; // @[OneHot.scala 32:28]
  wire [3:0] r_size = {_r_size_T_5,_r_size_T_7,_r_size_T_9,_r_size_T_10[1]}; // @[Cat.scala 33:92]
  reg [2:0] r_count_0; // @[ToTL.scala 102:28]
  reg [2:0] r_count_1; // @[ToTL.scala 102:28]
  wire [2:0] _GEN_1 = auto_in_ar_bits_id ? r_count_1 : r_count_0; // @[ToTL.scala 106:{50,50}]
  wire [3:0] r_id = {auto_in_ar_bits_id,_GEN_1[1:0],1'h0}; // @[Cat.scala 33:92]
  wire [29:0] _T_2 = 30'h7fff << r_size; // @[package.scala 235:71]
  wire [14:0] _T_4 = ~_T_2[14:0]; // @[package.scala 235:46]
  wire  _T_8 = ~reset; // @[ToTL.scala 109:14]
  wire [1:0] r_sel = 2'h1 << auto_in_ar_bits_id; // @[OneHot.scala 64:12]
  reg [7:0] beatsLeft; // @[Arbiter.scala 88:30]
  wire  idle = beatsLeft == 8'h0; // @[Arbiter.scala 89:28]
  wire  w_out_valid = auto_in_aw_valid & auto_in_w_valid; // @[ToTL.scala 146:34]
  wire [1:0] readys_valid = {w_out_valid,auto_in_ar_valid}; // @[Cat.scala 33:92]
  reg [1:0] readys_mask; // @[Arbiter.scala 24:23]
  wire [1:0] _readys_filter_T = ~readys_mask; // @[Arbiter.scala 25:30]
  wire [1:0] _readys_filter_T_1 = readys_valid & _readys_filter_T; // @[Arbiter.scala 25:28]
  wire [3:0] readys_filter = {_readys_filter_T_1,w_out_valid,auto_in_ar_valid}; // @[Cat.scala 33:92]
  wire [3:0] _GEN_16 = {{1'd0}, readys_filter[3:1]}; // @[package.scala 254:43]
  wire [3:0] _readys_unready_T_1 = readys_filter | _GEN_16; // @[package.scala 254:43]
  wire [3:0] _readys_unready_T_4 = {readys_mask, 2'h0}; // @[Arbiter.scala 26:66]
  wire [3:0] _GEN_17 = {{1'd0}, _readys_unready_T_1[3:1]}; // @[Arbiter.scala 26:58]
  wire [3:0] readys_unready = _GEN_17 | _readys_unready_T_4; // @[Arbiter.scala 26:58]
  wire [1:0] _readys_readys_T_2 = readys_unready[3:2] & readys_unready[1:0]; // @[Arbiter.scala 27:39]
  wire [1:0] readys_readys = ~_readys_readys_T_2; // @[Arbiter.scala 27:18]
  wire  readys_0 = readys_readys[0]; // @[Arbiter.scala 96:86]
  reg  state_0; // @[Arbiter.scala 117:26]
  wire  allowed_0 = idle ? readys_0 : state_0; // @[Arbiter.scala 122:24]
  wire  out_ready = auto_out_a_ready & allowed_0; // @[Arbiter.scala 124:31]
  wire  _T_12 = out_ready & auto_in_ar_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _r_count_0_T_1 = r_count_0 + 3'h1; // @[ToTL.scala 127:41]
  wire [2:0] _r_count_1_T_1 = r_count_1 + 3'h1; // @[ToTL.scala 127:41]
  wire [22:0] _w_size1_T_1 = 23'hff << auto_in_aw_bits_size; // @[Bundles.scala 33:21]
  wire [14:0] w_size1 = _w_size1_T_1[22:8]; // @[Bundles.scala 33:30]
  wire [15:0] _w_size_T = {w_size1, 1'h0}; // @[package.scala 233:35]
  wire [15:0] _w_size_T_1 = _w_size_T | 16'h1; // @[package.scala 233:40]
  wire [15:0] _w_size_T_2 = {1'h0,w_size1}; // @[Cat.scala 33:92]
  wire [15:0] _w_size_T_3 = ~_w_size_T_2; // @[package.scala 233:49]
  wire [15:0] _w_size_T_4 = _w_size_T_1 & _w_size_T_3; // @[package.scala 233:47]
  wire [7:0] w_size_hi = _w_size_T_4[15:8]; // @[OneHot.scala 30:18]
  wire [7:0] w_size_lo = _w_size_T_4[7:0]; // @[OneHot.scala 31:18]
  wire  _w_size_T_5 = |w_size_hi; // @[OneHot.scala 32:14]
  wire [7:0] _w_size_T_6 = w_size_hi | w_size_lo; // @[OneHot.scala 32:28]
  wire [3:0] w_size_hi_1 = _w_size_T_6[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] w_size_lo_1 = _w_size_T_6[3:0]; // @[OneHot.scala 31:18]
  wire  _w_size_T_7 = |w_size_hi_1; // @[OneHot.scala 32:14]
  wire [3:0] _w_size_T_8 = w_size_hi_1 | w_size_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] w_size_hi_2 = _w_size_T_8[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] w_size_lo_2 = _w_size_T_8[1:0]; // @[OneHot.scala 31:18]
  wire  _w_size_T_9 = |w_size_hi_2; // @[OneHot.scala 32:14]
  wire [1:0] _w_size_T_10 = w_size_hi_2 | w_size_lo_2; // @[OneHot.scala 32:28]
  wire [3:0] w_size = {_w_size_T_5,_w_size_T_7,_w_size_T_9,_w_size_T_10[1]}; // @[Cat.scala 33:92]
  reg [2:0] w_count_0; // @[ToTL.scala 135:28]
  reg [2:0] w_count_1; // @[ToTL.scala 135:28]
  wire [2:0] _GEN_5 = auto_in_aw_bits_id ? w_count_1 : w_count_0; // @[ToTL.scala 139:{50,50}]
  wire [3:0] w_id = {auto_in_aw_bits_id,_GEN_5[1:0],1'h1}; // @[Cat.scala 33:92]
  wire [29:0] _T_18 = 30'h7fff << w_size; // @[package.scala 235:71]
  wire [14:0] _T_20 = ~_T_18[14:0]; // @[package.scala 235:46]
  wire  readys_1 = readys_readys[1]; // @[Arbiter.scala 96:86]
  reg  state_1; // @[Arbiter.scala 117:26]
  wire  allowed_1 = idle ? readys_1 : state_1; // @[Arbiter.scala 122:24]
  wire  out_1_ready = auto_out_a_ready & allowed_1; // @[Arbiter.scala 124:31]
  wire  bundleIn_0_aw_ready = out_1_ready & auto_in_w_valid & auto_in_w_bits_last; // @[ToTL.scala 144:48]
  wire [1:0] w_sel = 2'h1 << auto_in_aw_bits_id; // @[OneHot.scala 64:12]
  wire  _T_36 = bundleIn_0_aw_ready & auto_in_aw_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _w_count_0_T_1 = w_count_0 + 3'h1; // @[ToTL.scala 163:41]
  wire [2:0] _w_count_1_T_1 = w_count_1 + 3'h1; // @[ToTL.scala 163:41]
  wire  latch = idle & auto_out_a_ready; // @[Arbiter.scala 90:24]
  wire [1:0] _readys_mask_T = readys_readys & readys_valid; // @[Arbiter.scala 29:29]
  wire [2:0] _readys_mask_T_1 = {_readys_mask_T, 1'h0}; // @[package.scala 245:48]
  wire [1:0] _readys_mask_T_3 = _readys_mask_T | _readys_mask_T_1[1:0]; // @[package.scala 245:43]
  wire  earlyWinner_0 = readys_0 & auto_in_ar_valid; // @[Arbiter.scala 98:79]
  wire  earlyWinner_1 = readys_1 & w_out_valid; // @[Arbiter.scala 98:79]
  wire  _prefixOR_T = earlyWinner_0 | earlyWinner_1; // @[Arbiter.scala 105:53]
  wire  _T_50 = auto_in_ar_valid | w_out_valid; // @[Arbiter.scala 108:36]
  wire  _T_51 = ~(auto_in_ar_valid | w_out_valid); // @[Arbiter.scala 108:15]
  wire  muxStateEarly_0 = idle ? earlyWinner_0 : state_0; // @[Arbiter.scala 118:30]
  wire  muxStateEarly_1 = idle ? earlyWinner_1 : state_1; // @[Arbiter.scala 118:30]
  wire  _sink_ACancel_earlyValid_T_3 = state_0 & auto_in_ar_valid | state_1 & w_out_valid; // @[Mux.scala 27:73]
  wire  sink_ACancel_earlyValid = idle ? _T_50 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 126:29]
  wire  _beatsLeft_T_2 = auto_out_a_ready & sink_ACancel_earlyValid; // @[ReadyValidCancel.scala 49:33]
  wire [7:0] _GEN_18 = {{7'd0}, _beatsLeft_T_2}; // @[Arbiter.scala 114:52]
  wire [7:0] _beatsLeft_T_4 = beatsLeft - _GEN_18; // @[Arbiter.scala 114:52]
  wire [15:0] _T_73 = muxStateEarly_0 ? auto_in_ar_bits_addr : 16'h0; // @[Mux.scala 27:73]
  wire [15:0] _T_74 = muxStateEarly_1 ? auto_in_aw_bits_addr : 16'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_76 = muxStateEarly_0 ? r_id : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_77 = muxStateEarly_1 ? w_id : 4'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_85 = muxStateEarly_0 ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_86 = muxStateEarly_1 ? 3'h1 : 3'h0; // @[Mux.scala 27:73]
  wire  d_hasData = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire  ok_r_ready = deq_io_enq_ready; // @[ToTL.scala 169:30 Decoupled.scala 379:17]
  wire  ok_b_ready = q_b_deq_io_enq_ready; // @[ToTL.scala 168:30 Decoupled.scala 379:17]
  reg [2:0] b_count_0; // @[ToTL.scala 197:28]
  reg [2:0] b_count_1; // @[ToTL.scala 197:28]
  wire  q_b_bits_id = q_b_deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  wire [2:0] _GEN_11 = q_b_bits_id ? b_count_1 : b_count_0; // @[ToTL.scala 198:{43,43}]
  wire [2:0] _GEN_13 = q_b_bits_id ? w_count_1 : w_count_0; // @[ToTL.scala 198:{43,43}]
  wire  b_allow = _GEN_11 != _GEN_13; // @[ToTL.scala 198:43]
  wire [1:0] b_sel = 2'h1 << q_b_bits_id; // @[OneHot.scala 64:12]
  wire  q_b_valid = q_b_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  wire  bundleIn_0_b_valid = q_b_valid & b_allow; // @[ToTL.scala 206:31]
  wire  _T_90 = auto_in_b_ready & bundleIn_0_b_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _b_count_0_T_1 = b_count_0 + 3'h1; // @[ToTL.scala 202:40]
  wire [2:0] _b_count_1_T_1 = b_count_1 + 3'h1; // @[ToTL.scala 202:40]
  Queue_171 deq ( // @[Decoupled.scala 375:21]
    .clock(deq_clock),
    .reset(deq_reset),
    .io_enq_ready(deq_io_enq_ready),
    .io_enq_valid(deq_io_enq_valid),
    .io_enq_bits_id(deq_io_enq_bits_id),
    .io_enq_bits_data(deq_io_enq_bits_data),
    .io_deq_ready(deq_io_deq_ready),
    .io_deq_valid(deq_io_deq_valid),
    .io_deq_bits_id(deq_io_deq_bits_id),
    .io_deq_bits_data(deq_io_deq_bits_data),
    .io_deq_bits_resp(deq_io_deq_bits_resp),
    .io_deq_bits_last(deq_io_deq_bits_last)
  );
  Queue_172 q_b_deq ( // @[Decoupled.scala 375:21]
    .clock(q_b_deq_clock),
    .reset(q_b_deq_reset),
    .io_enq_ready(q_b_deq_io_enq_ready),
    .io_enq_valid(q_b_deq_io_enq_valid),
    .io_enq_bits_id(q_b_deq_io_enq_bits_id),
    .io_deq_ready(q_b_deq_io_deq_ready),
    .io_deq_valid(q_b_deq_io_deq_valid),
    .io_deq_bits_id(q_b_deq_io_deq_bits_id),
    .io_deq_bits_resp(q_b_deq_io_deq_bits_resp)
  );
  assign auto_in_aw_ready = out_1_ready & auto_in_w_valid & auto_in_w_bits_last; // @[ToTL.scala 144:48]
  assign auto_in_w_ready = out_1_ready & auto_in_aw_valid; // @[ToTL.scala 145:34]
  assign auto_in_b_valid = q_b_valid & b_allow; // @[ToTL.scala 206:31]
  assign auto_in_b_bits_id = q_b_deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_b_bits_resp = q_b_deq_io_deq_bits_resp; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_ar_ready = auto_out_a_ready & allowed_0; // @[Arbiter.scala 124:31]
  assign auto_in_r_valid = deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_in_r_bits_id = deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_r_bits_data = deq_io_deq_bits_data; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_r_bits_resp = deq_io_deq_bits_resp; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_r_bits_last = deq_io_deq_bits_last; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_a_valid = idle ? _T_50 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 126:29]
  assign auto_out_a_bits_opcode = _T_85 | _T_86; // @[Mux.scala 27:73]
  assign auto_out_a_bits_source = _T_76 | _T_77; // @[Mux.scala 27:73]
  assign auto_out_a_bits_address = _T_73 | _T_74; // @[Mux.scala 27:73]
  assign auto_out_a_bits_data = muxStateEarly_1 ? auto_in_w_bits_data : 32'h0; // @[Mux.scala 27:73]
  assign auto_out_d_ready = d_hasData ? ok_r_ready : ok_b_ready; // @[ToTL.scala 175:25]
  assign deq_clock = clock;
  assign deq_reset = reset;
  assign deq_io_enq_valid = auto_out_d_valid & d_hasData; // @[ToTL.scala 176:33]
  assign deq_io_enq_bits_id = auto_out_d_bits_source[3]; // @[ToTL.scala 179:43]
  assign deq_io_enq_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign deq_io_deq_ready = auto_in_r_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign q_b_deq_clock = clock;
  assign q_b_deq_reset = reset;
  assign q_b_deq_io_enq_valid = auto_out_d_valid & ~d_hasData; // @[ToTL.scala 177:33]
  assign q_b_deq_io_enq_bits_id = auto_out_d_bits_source[3]; // @[ToTL.scala 188:43]
  assign q_b_deq_io_deq_ready = auto_in_b_ready & b_allow; // @[ToTL.scala 207:31]
  always @(posedge clock) begin
    if (reset) begin // @[ToTL.scala 102:28]
      r_count_0 <= 3'h0; // @[ToTL.scala 102:28]
    end else if (_T_12 & r_sel[0]) begin // @[ToTL.scala 127:32]
      r_count_0 <= _r_count_0_T_1; // @[ToTL.scala 127:36]
    end
    if (reset) begin // @[ToTL.scala 102:28]
      r_count_1 <= 3'h0; // @[ToTL.scala 102:28]
    end else if (_T_12 & r_sel[1]) begin // @[ToTL.scala 127:32]
      r_count_1 <= _r_count_1_T_1; // @[ToTL.scala 127:36]
    end
    if (reset) begin // @[Arbiter.scala 88:30]
      beatsLeft <= 8'h0; // @[Arbiter.scala 88:30]
    end else if (latch) begin // @[Arbiter.scala 114:23]
      beatsLeft <= 8'h0;
    end else begin
      beatsLeft <= _beatsLeft_T_4;
    end
    if (reset) begin // @[Arbiter.scala 24:23]
      readys_mask <= 2'h3; // @[Arbiter.scala 24:23]
    end else if (latch & |readys_valid) begin // @[Arbiter.scala 28:32]
      readys_mask <= _readys_mask_T_3; // @[Arbiter.scala 29:12]
    end
    if (reset) begin // @[Arbiter.scala 117:26]
      state_0 <= 1'h0; // @[Arbiter.scala 117:26]
    end else if (idle) begin // @[Arbiter.scala 118:30]
      state_0 <= earlyWinner_0;
    end
    if (reset) begin // @[ToTL.scala 135:28]
      w_count_0 <= 3'h0; // @[ToTL.scala 135:28]
    end else if (_T_36 & w_sel[0]) begin // @[ToTL.scala 163:32]
      w_count_0 <= _w_count_0_T_1; // @[ToTL.scala 163:36]
    end
    if (reset) begin // @[ToTL.scala 135:28]
      w_count_1 <= 3'h0; // @[ToTL.scala 135:28]
    end else if (_T_36 & w_sel[1]) begin // @[ToTL.scala 163:32]
      w_count_1 <= _w_count_1_T_1; // @[ToTL.scala 163:36]
    end
    if (reset) begin // @[Arbiter.scala 117:26]
      state_1 <= 1'h0; // @[Arbiter.scala 117:26]
    end else if (idle) begin // @[Arbiter.scala 118:30]
      state_1 <= earlyWinner_1;
    end
    if (reset) begin // @[ToTL.scala 197:28]
      b_count_0 <= 3'h0; // @[ToTL.scala 197:28]
    end else if (_T_90 & b_sel[0]) begin // @[ToTL.scala 202:31]
      b_count_0 <= _b_count_0_T_1; // @[ToTL.scala 202:35]
    end
    if (reset) begin // @[ToTL.scala 197:28]
      b_count_1 <= 3'h0; // @[ToTL.scala 197:28]
    end else if (_T_90 & b_sel[1]) begin // @[ToTL.scala 202:31]
      b_count_1 <= _b_count_1_T_1; // @[ToTL.scala 202:35]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~auto_in_ar_valid | r_size1 == _T_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToTL.scala:109 assert (!in.ar.valid || r_size1 === UIntToOH1(r_size, beatCountBits)) // because aligned\n"
            ); // @[ToTL.scala 109:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~auto_in_ar_valid | r_size1 == _T_4) & ~reset) begin
          $fatal; // @[ToTL.scala 109:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & ~(~auto_in_aw_valid | w_size1 == _T_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToTL.scala:142 assert (!in.aw.valid || w_size1 === UIntToOH1(w_size, beatCountBits)) // because aligned\n"
            ); // @[ToTL.scala 142:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~auto_in_aw_valid | w_size1 == _T_20) & _T_8) begin
          $fatal; // @[ToTL.scala 142:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & ~(~earlyWinner_0 | ~earlyWinner_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:106 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[Arbiter.scala 106:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~earlyWinner_0 | ~earlyWinner_1) & _T_8) begin
          $fatal; // @[Arbiter.scala 106:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & ~(~(auto_in_ar_valid | w_out_valid) | _prefixOR_T)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:108 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"
            ); // @[Arbiter.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(auto_in_ar_valid | w_out_valid) | _prefixOR_T) & _T_8) begin
          $fatal; // @[Arbiter.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & ~(_T_51 | _T_50)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:109 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"
            ); // @[Arbiter.scala 109:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_51 | _T_50) & _T_8) begin
          $fatal; // @[Arbiter.scala 109:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_173(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [14:0] io_enq_bits_extra_id,
  input         io_enq_bits_real_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [14:0] io_deq_bits_extra_id,
  output        io_deq_bits_real_last
);
  reg [14:0] ram_extra_id [0:3]; // @[Decoupled.scala 273:95]
  wire  ram_extra_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_extra_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [14:0] ram_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [14:0] ram_extra_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_extra_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_extra_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_extra_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_real_last [0:3]; // @[Decoupled.scala 273:95]
  wire  ram_real_last_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_real_last_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_real_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_real_last_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_real_last_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_real_last_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_real_last_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire  _GEN_13 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 318:26 280:27 318:35]
  wire  do_enq = empty ? _GEN_13 : _do_enq_T; // @[Decoupled.scala 315:17 280:27]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 315:17 317:14 281:27]
  assign ram_extra_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_extra_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_extra_id_io_deq_bits_MPORT_data = ram_extra_id[ram_extra_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_extra_id_MPORT_data = io_enq_bits_extra_id;
  assign ram_extra_id_MPORT_addr = enq_ptr_value;
  assign ram_extra_id_MPORT_mask = 1'h1;
  assign ram_extra_id_MPORT_en = empty ? _GEN_13 : _do_enq_T;
  assign ram_real_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_real_last_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_real_last_io_deq_bits_MPORT_data = ram_real_last[ram_real_last_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_real_last_MPORT_data = io_enq_bits_real_last;
  assign ram_real_last_MPORT_addr = enq_ptr_value;
  assign ram_real_last_MPORT_mask = 1'h1;
  assign ram_real_last_MPORT_en = empty ? _GEN_13 : _do_enq_T;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 302:16 314:{24,39}]
  assign io_deq_bits_extra_id = empty ? io_enq_bits_extra_id : ram_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_real_last = empty ? io_enq_bits_real_last : ram_real_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  always @(posedge clock) begin
    if (ram_extra_id_MPORT_en & ram_extra_id_MPORT_mask) begin
      ram_extra_id[ram_extra_id_MPORT_addr] <= ram_extra_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_real_last_MPORT_en & ram_real_last_MPORT_mask) begin
      ram_real_last[ram_real_last_MPORT_addr] <= ram_real_last_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      if (empty) begin // @[Decoupled.scala 315:17]
        if (io_deq_ready) begin // @[Decoupled.scala 318:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 318:35]
        end else begin
          maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
        end
      end else begin
        maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
      end
    end
  end
endmodule
module AXI4UserYanker_1(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [15:0] auto_in_aw_bits_addr,
  input  [2:0]  auto_in_aw_bits_size,
  input  [14:0] auto_in_aw_bits_echo_extra_id,
  input         auto_in_aw_bits_echo_real_last,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output        auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output [14:0] auto_in_b_bits_echo_extra_id,
  output        auto_in_b_bits_echo_real_last,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [15:0] auto_in_ar_bits_addr,
  input  [2:0]  auto_in_ar_bits_size,
  input  [14:0] auto_in_ar_bits_echo_extra_id,
  input         auto_in_ar_bits_echo_real_last,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output        auto_in_r_bits_id,
  output [31:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output [14:0] auto_in_r_bits_echo_extra_id,
  output        auto_in_r_bits_echo_real_last,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output        auto_out_aw_bits_id,
  output [15:0] auto_out_aw_bits_addr,
  output [2:0]  auto_out_aw_bits_size,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [31:0] auto_out_w_bits_data,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input         auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output        auto_out_ar_bits_id,
  output [15:0] auto_out_ar_bits_addr,
  output [2:0]  auto_out_ar_bits_size,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input         auto_out_r_bits_id,
  input  [31:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input         auto_out_r_bits_last
);
  wire  Queue_clock; // @[UserYanker.scala 50:17]
  wire  Queue_reset; // @[UserYanker.scala 50:17]
  wire  Queue_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [14:0] Queue_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_io_enq_bits_real_last; // @[UserYanker.scala 50:17]
  wire  Queue_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [14:0] Queue_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_io_deq_bits_real_last; // @[UserYanker.scala 50:17]
  wire  Queue_1_clock; // @[UserYanker.scala 50:17]
  wire  Queue_1_reset; // @[UserYanker.scala 50:17]
  wire  Queue_1_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_1_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [14:0] Queue_1_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_1_io_enq_bits_real_last; // @[UserYanker.scala 50:17]
  wire  Queue_1_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_1_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [14:0] Queue_1_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_1_io_deq_bits_real_last; // @[UserYanker.scala 50:17]
  wire  Queue_2_clock; // @[UserYanker.scala 50:17]
  wire  Queue_2_reset; // @[UserYanker.scala 50:17]
  wire  Queue_2_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_2_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [14:0] Queue_2_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_2_io_enq_bits_real_last; // @[UserYanker.scala 50:17]
  wire  Queue_2_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_2_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [14:0] Queue_2_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_2_io_deq_bits_real_last; // @[UserYanker.scala 50:17]
  wire  Queue_3_clock; // @[UserYanker.scala 50:17]
  wire  Queue_3_reset; // @[UserYanker.scala 50:17]
  wire  Queue_3_io_enq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_3_io_enq_valid; // @[UserYanker.scala 50:17]
  wire [14:0] Queue_3_io_enq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_3_io_enq_bits_real_last; // @[UserYanker.scala 50:17]
  wire  Queue_3_io_deq_ready; // @[UserYanker.scala 50:17]
  wire  Queue_3_io_deq_valid; // @[UserYanker.scala 50:17]
  wire [14:0] Queue_3_io_deq_bits_extra_id; // @[UserYanker.scala 50:17]
  wire  Queue_3_io_deq_bits_real_last; // @[UserYanker.scala 50:17]
  wire  _ar_ready_WIRE_0 = Queue_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _ar_ready_WIRE_1 = Queue_1_io_enq_ready; // @[UserYanker.scala 58:{29,29}]
  wire  _GEN_1 = auto_in_ar_bits_id ? _ar_ready_WIRE_1 : _ar_ready_WIRE_0; // @[UserYanker.scala 59:{36,36}]
  wire  _r_valid_WIRE_0 = Queue_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _r_valid_WIRE_1 = Queue_1_io_deq_valid; // @[UserYanker.scala 64:{28,28}]
  wire  _GEN_3 = auto_out_r_bits_id ? _r_valid_WIRE_1 : _r_valid_WIRE_0; // @[UserYanker.scala 66:{28,28}]
  wire  _T_3 = ~reset; // @[UserYanker.scala 66:14]
  wire  _r_bits_WIRE_0_real_last = Queue_io_deq_bits_real_last; // @[UserYanker.scala 65:{27,27}]
  wire  _r_bits_WIRE_1_real_last = Queue_1_io_deq_bits_real_last; // @[UserYanker.scala 65:{27,27}]
  wire [14:0] _r_bits_WIRE_0_extra_id = Queue_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [14:0] _r_bits_WIRE_1_extra_id = Queue_1_io_deq_bits_extra_id; // @[UserYanker.scala 65:{27,27}]
  wire [1:0] _arsel_T = 2'h1 << auto_in_ar_bits_id; // @[OneHot.scala 64:12]
  wire  arsel_0 = _arsel_T[0]; // @[UserYanker.scala 70:55]
  wire  arsel_1 = _arsel_T[1]; // @[UserYanker.scala 70:55]
  wire [1:0] _rsel_T = 2'h1 << auto_out_r_bits_id; // @[OneHot.scala 64:12]
  wire  rsel_0 = _rsel_T[0]; // @[UserYanker.scala 71:55]
  wire  rsel_1 = _rsel_T[1]; // @[UserYanker.scala 71:55]
  wire  _aw_ready_WIRE_0 = Queue_2_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _aw_ready_WIRE_1 = Queue_3_io_enq_ready; // @[UserYanker.scala 79:{29,29}]
  wire  _GEN_9 = auto_in_aw_bits_id ? _aw_ready_WIRE_1 : _aw_ready_WIRE_0; // @[UserYanker.scala 80:{36,36}]
  wire  _b_valid_WIRE_0 = Queue_2_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _b_valid_WIRE_1 = Queue_3_io_deq_valid; // @[UserYanker.scala 85:{28,28}]
  wire  _GEN_11 = auto_out_b_bits_id ? _b_valid_WIRE_1 : _b_valid_WIRE_0; // @[UserYanker.scala 87:{28,28}]
  wire  _b_bits_WIRE_0_real_last = Queue_2_io_deq_bits_real_last; // @[UserYanker.scala 86:{27,27}]
  wire  _b_bits_WIRE_1_real_last = Queue_3_io_deq_bits_real_last; // @[UserYanker.scala 86:{27,27}]
  wire [14:0] _b_bits_WIRE_0_extra_id = Queue_2_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [14:0] _b_bits_WIRE_1_extra_id = Queue_3_io_deq_bits_extra_id; // @[UserYanker.scala 86:{27,27}]
  wire [1:0] _awsel_T = 2'h1 << auto_in_aw_bits_id; // @[OneHot.scala 64:12]
  wire  awsel_0 = _awsel_T[0]; // @[UserYanker.scala 91:55]
  wire  awsel_1 = _awsel_T[1]; // @[UserYanker.scala 91:55]
  wire [1:0] _bsel_T = 2'h1 << auto_out_b_bits_id; // @[OneHot.scala 64:12]
  wire  bsel_0 = _bsel_T[0]; // @[UserYanker.scala 92:55]
  wire  bsel_1 = _bsel_T[1]; // @[UserYanker.scala 92:55]
  Queue_173 Queue ( // @[UserYanker.scala 50:17]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_extra_id(Queue_io_enq_bits_extra_id),
    .io_enq_bits_real_last(Queue_io_enq_bits_real_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_extra_id(Queue_io_deq_bits_extra_id),
    .io_deq_bits_real_last(Queue_io_deq_bits_real_last)
  );
  Queue_173 Queue_1 ( // @[UserYanker.scala 50:17]
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_extra_id(Queue_1_io_enq_bits_extra_id),
    .io_enq_bits_real_last(Queue_1_io_enq_bits_real_last),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_extra_id(Queue_1_io_deq_bits_extra_id),
    .io_deq_bits_real_last(Queue_1_io_deq_bits_real_last)
  );
  Queue_173 Queue_2 ( // @[UserYanker.scala 50:17]
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_extra_id(Queue_2_io_enq_bits_extra_id),
    .io_enq_bits_real_last(Queue_2_io_enq_bits_real_last),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_extra_id(Queue_2_io_deq_bits_extra_id),
    .io_deq_bits_real_last(Queue_2_io_deq_bits_real_last)
  );
  Queue_173 Queue_3 ( // @[UserYanker.scala 50:17]
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits_extra_id(Queue_3_io_enq_bits_extra_id),
    .io_enq_bits_real_last(Queue_3_io_enq_bits_real_last),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits_extra_id(Queue_3_io_deq_bits_extra_id),
    .io_deq_bits_real_last(Queue_3_io_deq_bits_real_last)
  );
  assign auto_in_aw_ready = auto_out_aw_ready & _GEN_9; // @[UserYanker.scala 80:36]
  assign auto_in_w_ready = auto_out_w_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_b_valid = auto_out_b_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_b_bits_id = auto_out_b_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_b_bits_echo_extra_id = auto_out_b_bits_id ? _b_bits_WIRE_1_extra_id : _b_bits_WIRE_0_extra_id; // @[BundleMap.scala 247:{19,19}]
  assign auto_in_b_bits_echo_real_last = auto_out_b_bits_id ? _b_bits_WIRE_1_real_last : _b_bits_WIRE_0_real_last; // @[BundleMap.scala 247:{19,19}]
  assign auto_in_ar_ready = auto_out_ar_ready & _GEN_1; // @[UserYanker.scala 59:36]
  assign auto_in_r_valid = auto_out_r_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_bits_id = auto_out_r_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_bits_echo_extra_id = auto_out_r_bits_id ? _r_bits_WIRE_1_extra_id : _r_bits_WIRE_0_extra_id; // @[BundleMap.scala 247:{19,19}]
  assign auto_in_r_bits_echo_real_last = auto_out_r_bits_id ? _r_bits_WIRE_1_real_last : _r_bits_WIRE_0_real_last; // @[BundleMap.scala 247:{19,19}]
  assign auto_in_r_bits_last = auto_out_r_bits_last; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_out_aw_valid = auto_in_aw_valid & _GEN_9; // @[UserYanker.scala 81:36]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_size = auto_in_aw_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_w_valid = auto_in_w_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_b_ready = auto_in_b_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_valid = auto_in_ar_valid & _GEN_1; // @[UserYanker.scala 60:36]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_r_ready = auto_in_r_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_0; // @[UserYanker.scala 74:53]
  assign Queue_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_io_enq_bits_real_last = auto_in_ar_bits_echo_real_last; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_0 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_1; // @[UserYanker.scala 74:53]
  assign Queue_1_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_1_io_enq_bits_real_last = auto_in_ar_bits_echo_real_last; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_1_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_1 & auto_out_r_bits_last; // @[UserYanker.scala 73:58]
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign Queue_2_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_0; // @[UserYanker.scala 95:53]
  assign Queue_2_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_2_io_enq_bits_real_last = auto_in_aw_bits_echo_real_last; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_2_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_0; // @[UserYanker.scala 94:53]
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign Queue_3_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_1; // @[UserYanker.scala 95:53]
  assign Queue_3_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_3_io_enq_bits_real_last = auto_in_aw_bits_echo_real_last; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign Queue_3_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_1; // @[UserYanker.scala 94:53]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~auto_out_r_valid | _GEN_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at UserYanker.scala:66 assert (!out.r.valid || r_valid) // Q must be ready faster than the response\n"
            ); // @[UserYanker.scala 66:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~auto_out_r_valid | _GEN_3) & ~reset) begin
          $fatal; // @[UserYanker.scala 66:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3 & ~(~auto_out_b_valid | _GEN_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at UserYanker.scala:87 assert (!out.b.valid || b_valid) // Q must be ready faster than the response\n"
            ); // @[UserYanker.scala 87:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~auto_out_b_valid | _GEN_11) & _T_3) begin
          $fatal; // @[UserYanker.scala 87:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_177(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_id,
  input  [15:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_len,
  input  [2:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_burst,
  input  [14:0] io_enq_bits_echo_extra_id,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_id,
  output [15:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_len,
  output [2:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_burst,
  output [14:0] io_deq_bits_echo_extra_id
);
  reg  ram_id [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [15:0] ram_addr [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_addr_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_addr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [15:0] ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [15:0] ram_addr_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_addr_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_addr_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_addr_MPORT_en; // @[Decoupled.scala 273:95]
  reg [7:0] ram_len [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_len_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_len_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [7:0] ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [7:0] ram_len_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_len_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_len_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_len_MPORT_en; // @[Decoupled.scala 273:95]
  reg [2:0] ram_size [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_size_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_burst [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_burst_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_burst_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_burst_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_burst_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_burst_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_burst_MPORT_en; // @[Decoupled.scala 273:95]
  reg [14:0] ram_echo_extra_id [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_echo_extra_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_echo_extra_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [14:0] ram_echo_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [14:0] ram_echo_extra_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_echo_extra_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_echo_extra_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_echo_extra_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 278:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_18 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 318:26 280:27 318:35]
  wire  do_enq = empty ? _GEN_18 : _do_enq_T; // @[Decoupled.scala 315:17 280:27]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 315:17 317:14 281:27]
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = 1'h0;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = empty ? _GEN_18 : _do_enq_T;
  assign ram_addr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_addr_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = 1'h0;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = empty ? _GEN_18 : _do_enq_T;
  assign ram_len_io_deq_bits_MPORT_en = 1'h1;
  assign ram_len_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_len_io_deq_bits_MPORT_data = ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_len_MPORT_data = io_enq_bits_len;
  assign ram_len_MPORT_addr = 1'h0;
  assign ram_len_MPORT_mask = 1'h1;
  assign ram_len_MPORT_en = empty ? _GEN_18 : _do_enq_T;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = 1'h0;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = empty ? _GEN_18 : _do_enq_T;
  assign ram_burst_io_deq_bits_MPORT_en = 1'h1;
  assign ram_burst_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_burst_io_deq_bits_MPORT_data = ram_burst[ram_burst_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_burst_MPORT_data = io_enq_bits_burst;
  assign ram_burst_MPORT_addr = 1'h0;
  assign ram_burst_MPORT_mask = 1'h1;
  assign ram_burst_MPORT_en = empty ? _GEN_18 : _do_enq_T;
  assign ram_echo_extra_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_echo_extra_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_echo_extra_id_io_deq_bits_MPORT_data = ram_echo_extra_id[ram_echo_extra_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_echo_extra_id_MPORT_data = io_enq_bits_echo_extra_id;
  assign ram_echo_extra_id_MPORT_addr = 1'h0;
  assign ram_echo_extra_id_MPORT_mask = 1'h1;
  assign ram_echo_extra_id_MPORT_en = empty ? _GEN_18 : _do_enq_T;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 302:16 314:{24,39}]
  assign io_deq_bits_id = empty ? io_enq_bits_id : ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_addr = empty ? io_enq_bits_addr : ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_len = empty ? io_enq_bits_len : ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_size = empty ? io_enq_bits_size : ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_burst = empty ? io_enq_bits_burst : ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_echo_extra_id = empty ? io_enq_bits_echo_extra_id : ram_echo_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_len_MPORT_en & ram_len_MPORT_mask) begin
      ram_len[ram_len_MPORT_addr] <= ram_len_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_burst_MPORT_en & ram_burst_MPORT_mask) begin
      ram_burst[ram_burst_MPORT_addr] <= ram_burst_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_echo_extra_id_MPORT_en & ram_echo_extra_id_MPORT_mask) begin
      ram_echo_extra_id[ram_echo_extra_id_MPORT_addr] <= ram_echo_extra_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      if (empty) begin // @[Decoupled.scala 315:17]
        if (io_deq_ready) begin // @[Decoupled.scala 318:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 318:35]
        end else begin
          maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
        end
      end else begin
        maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
      end
    end
  end
endmodule
module Queue_179(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] ram_data [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [31:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [31:0] ram_data_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_last [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_en; // @[Decoupled.scala 273:95]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 278:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_11 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 318:26 280:27 318:35]
  wire  do_enq = empty ? _GEN_11 : _do_enq_T; // @[Decoupled.scala 315:17 280:27]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 315:17 317:14 281:27]
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = 1'h0;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = empty ? _GEN_11 : _do_enq_T;
  assign ram_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_last_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_last_io_deq_bits_MPORT_data = ram_last[ram_last_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_last_MPORT_data = io_enq_bits_last;
  assign ram_last_MPORT_addr = 1'h0;
  assign ram_last_MPORT_mask = 1'h1;
  assign ram_last_MPORT_en = empty ? _GEN_11 : _do_enq_T;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 302:16 314:{24,39}]
  assign io_deq_bits_data = empty ? io_enq_bits_data : ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_last = empty ? io_enq_bits_last : ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  always @(posedge clock) begin
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_last_MPORT_en & ram_last_MPORT_mask) begin
      ram_last[ram_last_MPORT_addr] <= ram_last_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      if (empty) begin // @[Decoupled.scala 315:17]
        if (io_deq_ready) begin // @[Decoupled.scala 318:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 318:35]
        end else begin
          maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
        end
      end else begin
        maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
      end
    end
  end
endmodule
module AXI4Fragmenter(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [15:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [1:0]  auto_in_aw_bits_burst,
  input  [14:0] auto_in_aw_bits_echo_extra_id,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output        auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output [14:0] auto_in_b_bits_echo_extra_id,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [15:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [1:0]  auto_in_ar_bits_burst,
  input  [14:0] auto_in_ar_bits_echo_extra_id,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output        auto_in_r_bits_id,
  output [31:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output [14:0] auto_in_r_bits_echo_extra_id,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output        auto_out_aw_bits_id,
  output [15:0] auto_out_aw_bits_addr,
  output [2:0]  auto_out_aw_bits_size,
  output [14:0] auto_out_aw_bits_echo_extra_id,
  output        auto_out_aw_bits_echo_real_last,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [31:0] auto_out_w_bits_data,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input         auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input  [14:0] auto_out_b_bits_echo_extra_id,
  input         auto_out_b_bits_echo_real_last,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output        auto_out_ar_bits_id,
  output [15:0] auto_out_ar_bits_addr,
  output [2:0]  auto_out_ar_bits_size,
  output [14:0] auto_out_ar_bits_echo_extra_id,
  output        auto_out_ar_bits_echo_real_last,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input         auto_out_r_bits_id,
  input  [31:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input  [14:0] auto_out_r_bits_echo_extra_id,
  input         auto_out_r_bits_echo_real_last,
  input         auto_out_r_bits_last
);
  wire  deq_clock; // @[Decoupled.scala 375:21]
  wire  deq_reset; // @[Decoupled.scala 375:21]
  wire  deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire  deq_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire [15:0] deq_io_enq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] deq_io_enq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] deq_io_enq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] deq_io_enq_bits_burst; // @[Decoupled.scala 375:21]
  wire [14:0] deq_io_enq_bits_echo_extra_id; // @[Decoupled.scala 375:21]
  wire  deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire  deq_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [15:0] deq_io_deq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] deq_io_deq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] deq_io_deq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] deq_io_deq_bits_burst; // @[Decoupled.scala 375:21]
  wire [14:0] deq_io_deq_bits_echo_extra_id; // @[Decoupled.scala 375:21]
  wire  deq_1_clock; // @[Decoupled.scala 375:21]
  wire  deq_1_reset; // @[Decoupled.scala 375:21]
  wire  deq_1_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  deq_1_io_enq_valid; // @[Decoupled.scala 375:21]
  wire  deq_1_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire [15:0] deq_1_io_enq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] deq_1_io_enq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] deq_1_io_enq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] deq_1_io_enq_bits_burst; // @[Decoupled.scala 375:21]
  wire [14:0] deq_1_io_enq_bits_echo_extra_id; // @[Decoupled.scala 375:21]
  wire  deq_1_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  deq_1_io_deq_valid; // @[Decoupled.scala 375:21]
  wire  deq_1_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [15:0] deq_1_io_deq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] deq_1_io_deq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] deq_1_io_deq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] deq_1_io_deq_bits_burst; // @[Decoupled.scala 375:21]
  wire [14:0] deq_1_io_deq_bits_echo_extra_id; // @[Decoupled.scala 375:21]
  wire  in_w_deq_clock; // @[Decoupled.scala 375:21]
  wire  in_w_deq_reset; // @[Decoupled.scala 375:21]
  wire  in_w_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  in_w_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [31:0] in_w_deq_io_enq_bits_data; // @[Decoupled.scala 375:21]
  wire  in_w_deq_io_enq_bits_last; // @[Decoupled.scala 375:21]
  wire  in_w_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  in_w_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [31:0] in_w_deq_io_deq_bits_data; // @[Decoupled.scala 375:21]
  wire  in_w_deq_io_deq_bits_last; // @[Decoupled.scala 375:21]
  reg  busy; // @[Fragmenter.scala 65:29]
  reg [15:0] r_addr; // @[Fragmenter.scala 66:25]
  reg [7:0] r_len; // @[Fragmenter.scala 67:25]
  wire [7:0] irr_bits_len = deq_io_deq_bits_len; // @[Decoupled.scala 414:19 415:14]
  wire [7:0] len = busy ? r_len : irr_bits_len; // @[Fragmenter.scala 69:23]
  wire [15:0] irr_bits_addr = deq_io_deq_bits_addr; // @[Decoupled.scala 414:19 415:14]
  wire [15:0] addr = busy ? r_addr : irr_bits_addr; // @[Fragmenter.scala 70:23]
  wire [1:0] irr_bits_burst = deq_io_deq_bits_burst; // @[Decoupled.scala 414:19 415:14]
  wire  fixed = irr_bits_burst == 2'h0; // @[Fragmenter.scala 97:34]
  wire [2:0] irr_bits_size = deq_io_deq_bits_size; // @[Decoupled.scala 414:19 415:14]
  wire [15:0] _inc_addr_T = 16'h1 << irr_bits_size; // @[Fragmenter.scala 105:38]
  wire [15:0] inc_addr = addr + _inc_addr_T; // @[Fragmenter.scala 105:29]
  wire [15:0] _wrapMask_T = {irr_bits_len,8'hff}; // @[Cat.scala 33:92]
  wire [22:0] _GEN_1 = {{7'd0}, _wrapMask_T}; // @[Bundles.scala 33:21]
  wire [22:0] _wrapMask_T_1 = _GEN_1 << irr_bits_size; // @[Bundles.scala 33:21]
  wire [14:0] wrapMask = _wrapMask_T_1[22:8]; // @[Bundles.scala 33:30]
  wire [15:0] _GEN_20 = {{1'd0}, wrapMask}; // @[Fragmenter.scala 109:33]
  wire [15:0] _mux_addr_T = inc_addr & _GEN_20; // @[Fragmenter.scala 109:33]
  wire [15:0] _mux_addr_T_1 = ~irr_bits_addr; // @[Fragmenter.scala 109:49]
  wire [15:0] _mux_addr_T_2 = _mux_addr_T_1 | _GEN_20; // @[Fragmenter.scala 109:62]
  wire [15:0] _mux_addr_T_3 = ~_mux_addr_T_2; // @[Fragmenter.scala 109:47]
  wire [15:0] _mux_addr_T_4 = _mux_addr_T | _mux_addr_T_3; // @[Fragmenter.scala 109:45]
  wire  ar_last = 8'h0 == len; // @[Fragmenter.scala 115:27]
  wire [15:0] _out_bits_addr_T = ~addr; // @[Fragmenter.scala 127:28]
  wire [8:0] _out_bits_addr_T_2 = 9'h3 << irr_bits_size; // @[package.scala 235:71]
  wire [1:0] _out_bits_addr_T_4 = ~_out_bits_addr_T_2[1:0]; // @[package.scala 235:46]
  wire [15:0] _GEN_22 = {{14'd0}, _out_bits_addr_T_4}; // @[Fragmenter.scala 127:34]
  wire [15:0] _out_bits_addr_T_5 = _out_bits_addr_T | _GEN_22; // @[Fragmenter.scala 127:34]
  wire  irr_valid = deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  wire  _T_2 = auto_out_ar_ready & irr_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _GEN_23 = {{1'd0}, len}; // @[Fragmenter.scala 132:25]
  wire [8:0] _r_len_T_1 = _GEN_23 - 9'h1; // @[Fragmenter.scala 132:25]
  wire [8:0] _GEN_4 = _T_2 ? _r_len_T_1 : {{1'd0}, r_len}; // @[Fragmenter.scala 129:25 132:18 67:25]
  reg  busy_1; // @[Fragmenter.scala 65:29]
  reg [15:0] r_addr_1; // @[Fragmenter.scala 66:25]
  reg [7:0] r_len_1; // @[Fragmenter.scala 67:25]
  wire [7:0] irr_1_bits_len = deq_1_io_deq_bits_len; // @[Decoupled.scala 414:19 415:14]
  wire [7:0] len_1 = busy_1 ? r_len_1 : irr_1_bits_len; // @[Fragmenter.scala 69:23]
  wire [15:0] irr_1_bits_addr = deq_1_io_deq_bits_addr; // @[Decoupled.scala 414:19 415:14]
  wire [15:0] addr_1 = busy_1 ? r_addr_1 : irr_1_bits_addr; // @[Fragmenter.scala 70:23]
  wire [1:0] irr_1_bits_burst = deq_1_io_deq_bits_burst; // @[Decoupled.scala 414:19 415:14]
  wire  fixed_1 = irr_1_bits_burst == 2'h0; // @[Fragmenter.scala 97:34]
  wire [2:0] irr_1_bits_size = deq_1_io_deq_bits_size; // @[Decoupled.scala 414:19 415:14]
  wire [15:0] _inc_addr_T_2 = 16'h1 << irr_1_bits_size; // @[Fragmenter.scala 105:38]
  wire [15:0] inc_addr_1 = addr_1 + _inc_addr_T_2; // @[Fragmenter.scala 105:29]
  wire [15:0] _wrapMask_T_2 = {irr_1_bits_len,8'hff}; // @[Cat.scala 33:92]
  wire [22:0] _GEN_3 = {{7'd0}, _wrapMask_T_2}; // @[Bundles.scala 33:21]
  wire [22:0] _wrapMask_T_3 = _GEN_3 << irr_1_bits_size; // @[Bundles.scala 33:21]
  wire [14:0] wrapMask_1 = _wrapMask_T_3[22:8]; // @[Bundles.scala 33:30]
  wire [15:0] _GEN_28 = {{1'd0}, wrapMask_1}; // @[Fragmenter.scala 109:33]
  wire [15:0] _mux_addr_T_5 = inc_addr_1 & _GEN_28; // @[Fragmenter.scala 109:33]
  wire [15:0] _mux_addr_T_6 = ~irr_1_bits_addr; // @[Fragmenter.scala 109:49]
  wire [15:0] _mux_addr_T_7 = _mux_addr_T_6 | _GEN_28; // @[Fragmenter.scala 109:62]
  wire [15:0] _mux_addr_T_8 = ~_mux_addr_T_7; // @[Fragmenter.scala 109:47]
  wire [15:0] _mux_addr_T_9 = _mux_addr_T_5 | _mux_addr_T_8; // @[Fragmenter.scala 109:45]
  wire  aw_last = 8'h0 == len_1; // @[Fragmenter.scala 115:27]
  reg [8:0] w_counter; // @[Fragmenter.scala 169:30]
  wire  w_idle = w_counter == 9'h0; // @[Fragmenter.scala 170:30]
  reg  wbeats_latched; // @[Fragmenter.scala 155:35]
  wire  _in_aw_ready_T = w_idle | wbeats_latched; // @[Fragmenter.scala 163:52]
  wire  in_aw_ready = auto_out_aw_ready & (w_idle | wbeats_latched); // @[Fragmenter.scala 163:35]
  wire [15:0] _out_bits_addr_T_7 = ~addr_1; // @[Fragmenter.scala 127:28]
  wire [8:0] _out_bits_addr_T_9 = 9'h3 << irr_1_bits_size; // @[package.scala 235:71]
  wire [1:0] _out_bits_addr_T_11 = ~_out_bits_addr_T_9[1:0]; // @[package.scala 235:46]
  wire [15:0] _GEN_30 = {{14'd0}, _out_bits_addr_T_11}; // @[Fragmenter.scala 127:34]
  wire [15:0] _out_bits_addr_T_12 = _out_bits_addr_T_7 | _GEN_30; // @[Fragmenter.scala 127:34]
  wire  irr_1_valid = deq_1_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  wire  _T_5 = in_aw_ready & irr_1_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _GEN_31 = {{1'd0}, len_1}; // @[Fragmenter.scala 132:25]
  wire [8:0] _r_len_T_3 = _GEN_31 - 9'h1; // @[Fragmenter.scala 132:25]
  wire [8:0] _GEN_9 = _T_5 ? _r_len_T_3 : {{1'd0}, r_len_1}; // @[Fragmenter.scala 129:25 132:18 67:25]
  wire  wbeats_valid = irr_1_valid & ~wbeats_latched; // @[Fragmenter.scala 164:35]
  wire  _GEN_10 = wbeats_valid & w_idle | wbeats_latched; // @[Fragmenter.scala 155:35 158:{43,60}]
  wire  x1_aw_valid = irr_1_valid & _in_aw_ready_T; // @[Fragmenter.scala 162:35]
  wire  _T_7 = auto_out_aw_ready & x1_aw_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _w_todo_T = wbeats_valid ? 9'h1 : 9'h0; // @[Fragmenter.scala 171:35]
  wire [8:0] w_todo = w_idle ? _w_todo_T : w_counter; // @[Fragmenter.scala 171:23]
  wire  w_last = w_todo == 9'h1; // @[Fragmenter.scala 172:27]
  wire  in_w_valid = in_w_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  wire  _x1_w_valid_T_1 = ~w_idle | wbeats_valid; // @[Fragmenter.scala 178:51]
  wire  x1_w_valid = in_w_valid & (~w_idle | wbeats_valid); // @[Fragmenter.scala 178:33]
  wire  _w_counter_T = auto_out_w_ready & x1_w_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _GEN_32 = {{8'd0}, _w_counter_T}; // @[Fragmenter.scala 173:27]
  wire [8:0] _w_counter_T_2 = w_todo - _GEN_32; // @[Fragmenter.scala 173:27]
  wire  _T_13 = ~reset; // @[Fragmenter.scala 174:14]
  wire  in_w_bits_last = in_w_deq_io_deq_bits_last; // @[Decoupled.scala 414:19 415:14]
  wire  x1_b_ready = auto_in_b_ready | ~auto_out_b_bits_echo_real_last; // @[Fragmenter.scala 194:33]
  reg [1:0] error_0; // @[Fragmenter.scala 197:26]
  reg [1:0] error_1; // @[Fragmenter.scala 197:26]
  wire [1:0] _GEN_13 = auto_out_b_bits_id ? error_1 : error_0; // @[Fragmenter.scala 198:{41,41}]
  wire [1:0] _T_22 = 2'h1 << auto_out_b_bits_id; // @[OneHot.scala 64:12]
  wire  _T_26 = x1_b_ready & auto_out_b_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _error_0_T = error_0 | auto_out_b_bits_resp; // @[Fragmenter.scala 200:64]
  wire [1:0] _error_1_T = error_1 | auto_out_b_bits_resp; // @[Fragmenter.scala 200:64]
  Queue_177 deq ( // @[Decoupled.scala 375:21]
    .clock(deq_clock),
    .reset(deq_reset),
    .io_enq_ready(deq_io_enq_ready),
    .io_enq_valid(deq_io_enq_valid),
    .io_enq_bits_id(deq_io_enq_bits_id),
    .io_enq_bits_addr(deq_io_enq_bits_addr),
    .io_enq_bits_len(deq_io_enq_bits_len),
    .io_enq_bits_size(deq_io_enq_bits_size),
    .io_enq_bits_burst(deq_io_enq_bits_burst),
    .io_enq_bits_echo_extra_id(deq_io_enq_bits_echo_extra_id),
    .io_deq_ready(deq_io_deq_ready),
    .io_deq_valid(deq_io_deq_valid),
    .io_deq_bits_id(deq_io_deq_bits_id),
    .io_deq_bits_addr(deq_io_deq_bits_addr),
    .io_deq_bits_len(deq_io_deq_bits_len),
    .io_deq_bits_size(deq_io_deq_bits_size),
    .io_deq_bits_burst(deq_io_deq_bits_burst),
    .io_deq_bits_echo_extra_id(deq_io_deq_bits_echo_extra_id)
  );
  Queue_177 deq_1 ( // @[Decoupled.scala 375:21]
    .clock(deq_1_clock),
    .reset(deq_1_reset),
    .io_enq_ready(deq_1_io_enq_ready),
    .io_enq_valid(deq_1_io_enq_valid),
    .io_enq_bits_id(deq_1_io_enq_bits_id),
    .io_enq_bits_addr(deq_1_io_enq_bits_addr),
    .io_enq_bits_len(deq_1_io_enq_bits_len),
    .io_enq_bits_size(deq_1_io_enq_bits_size),
    .io_enq_bits_burst(deq_1_io_enq_bits_burst),
    .io_enq_bits_echo_extra_id(deq_1_io_enq_bits_echo_extra_id),
    .io_deq_ready(deq_1_io_deq_ready),
    .io_deq_valid(deq_1_io_deq_valid),
    .io_deq_bits_id(deq_1_io_deq_bits_id),
    .io_deq_bits_addr(deq_1_io_deq_bits_addr),
    .io_deq_bits_len(deq_1_io_deq_bits_len),
    .io_deq_bits_size(deq_1_io_deq_bits_size),
    .io_deq_bits_burst(deq_1_io_deq_bits_burst),
    .io_deq_bits_echo_extra_id(deq_1_io_deq_bits_echo_extra_id)
  );
  Queue_179 in_w_deq ( // @[Decoupled.scala 375:21]
    .clock(in_w_deq_clock),
    .reset(in_w_deq_reset),
    .io_enq_ready(in_w_deq_io_enq_ready),
    .io_enq_valid(in_w_deq_io_enq_valid),
    .io_enq_bits_data(in_w_deq_io_enq_bits_data),
    .io_enq_bits_last(in_w_deq_io_enq_bits_last),
    .io_deq_ready(in_w_deq_io_deq_ready),
    .io_deq_valid(in_w_deq_io_deq_valid),
    .io_deq_bits_data(in_w_deq_io_deq_bits_data),
    .io_deq_bits_last(in_w_deq_io_deq_bits_last)
  );
  assign auto_in_aw_ready = deq_1_io_enq_ready; // @[Nodes.scala 1215:84 Decoupled.scala 379:17]
  assign auto_in_w_ready = in_w_deq_io_enq_ready; // @[Nodes.scala 1215:84 Decoupled.scala 379:17]
  assign auto_in_b_valid = auto_out_b_valid & auto_out_b_bits_echo_real_last; // @[Fragmenter.scala 193:33]
  assign auto_in_b_bits_id = auto_out_b_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp | _GEN_13; // @[Fragmenter.scala 198:41]
  assign auto_in_b_bits_echo_extra_id = auto_out_b_bits_echo_extra_id; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_ar_ready = deq_io_enq_ready; // @[Nodes.scala 1215:84 Decoupled.scala 379:17]
  assign auto_in_r_valid = auto_out_r_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_bits_id = auto_out_r_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_bits_echo_extra_id = auto_out_r_bits_echo_extra_id; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_bits_last = auto_out_r_bits_last & auto_out_r_bits_echo_real_last; // @[Fragmenter.scala 188:41]
  assign auto_out_aw_valid = irr_1_valid & _in_aw_ready_T; // @[Fragmenter.scala 162:35]
  assign auto_out_aw_bits_id = deq_1_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_addr = ~_out_bits_addr_T_12; // @[Fragmenter.scala 127:26]
  assign auto_out_aw_bits_size = deq_1_io_deq_bits_size; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_echo_extra_id = deq_1_io_deq_bits_echo_extra_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_echo_real_last = 8'h0 == len_1; // @[Fragmenter.scala 115:27]
  assign auto_out_w_valid = in_w_valid & (~w_idle | wbeats_valid); // @[Fragmenter.scala 178:33]
  assign auto_out_w_bits_data = in_w_deq_io_deq_bits_data; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_w_bits_last = w_todo == 9'h1; // @[Fragmenter.scala 172:27]
  assign auto_out_b_ready = auto_in_b_ready | ~auto_out_b_bits_echo_real_last; // @[Fragmenter.scala 194:33]
  assign auto_out_ar_valid = deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_out_ar_bits_id = deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_addr = ~_out_bits_addr_T_5; // @[Fragmenter.scala 127:26]
  assign auto_out_ar_bits_size = deq_io_deq_bits_size; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_echo_extra_id = deq_io_deq_bits_echo_extra_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_echo_real_last = 8'h0 == len; // @[Fragmenter.scala 115:27]
  assign auto_out_r_ready = auto_in_r_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign deq_clock = clock;
  assign deq_reset = reset;
  assign deq_io_enq_valid = auto_in_ar_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign deq_io_enq_bits_id = auto_in_ar_bits_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign deq_io_enq_bits_addr = auto_in_ar_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign deq_io_enq_bits_len = auto_in_ar_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign deq_io_enq_bits_size = auto_in_ar_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign deq_io_enq_bits_burst = auto_in_ar_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign deq_io_enq_bits_echo_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign deq_io_deq_ready = auto_out_ar_ready & ar_last; // @[Fragmenter.scala 116:30]
  assign deq_1_clock = clock;
  assign deq_1_reset = reset;
  assign deq_1_io_enq_valid = auto_in_aw_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign deq_1_io_enq_bits_id = auto_in_aw_bits_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign deq_1_io_enq_bits_addr = auto_in_aw_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign deq_1_io_enq_bits_len = auto_in_aw_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign deq_1_io_enq_bits_size = auto_in_aw_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign deq_1_io_enq_bits_burst = auto_in_aw_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign deq_1_io_enq_bits_echo_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign deq_1_io_deq_ready = in_aw_ready & aw_last; // @[Fragmenter.scala 116:30]
  assign in_w_deq_clock = clock;
  assign in_w_deq_reset = reset;
  assign in_w_deq_io_enq_valid = auto_in_w_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign in_w_deq_io_enq_bits_data = auto_in_w_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign in_w_deq_io_enq_bits_last = auto_in_w_bits_last; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign in_w_deq_io_deq_ready = auto_out_w_ready & _x1_w_valid_T_1; // @[Fragmenter.scala 179:33]
  always @(posedge clock) begin
    if (reset) begin // @[Fragmenter.scala 65:29]
      busy <= 1'h0; // @[Fragmenter.scala 65:29]
    end else if (_T_2) begin // @[Fragmenter.scala 129:25]
      busy <= ~ar_last; // @[Fragmenter.scala 130:16]
    end
    if (_T_2) begin // @[Fragmenter.scala 129:25]
      if (fixed) begin // @[Fragmenter.scala 111:60]
        r_addr <= irr_bits_addr; // @[Fragmenter.scala 112:20]
      end else if (irr_bits_burst == 2'h2) begin // @[Fragmenter.scala 108:59]
        r_addr <= _mux_addr_T_4; // @[Fragmenter.scala 109:20]
      end else begin
        r_addr <= inc_addr; // @[Fragmenter.scala 107:35]
      end
    end
    r_len <= _GEN_4[7:0];
    if (reset) begin // @[Fragmenter.scala 65:29]
      busy_1 <= 1'h0; // @[Fragmenter.scala 65:29]
    end else if (_T_5) begin // @[Fragmenter.scala 129:25]
      busy_1 <= ~aw_last; // @[Fragmenter.scala 130:16]
    end
    if (_T_5) begin // @[Fragmenter.scala 129:25]
      if (fixed_1) begin // @[Fragmenter.scala 111:60]
        r_addr_1 <= irr_1_bits_addr; // @[Fragmenter.scala 112:20]
      end else if (irr_1_bits_burst == 2'h2) begin // @[Fragmenter.scala 108:59]
        r_addr_1 <= _mux_addr_T_9; // @[Fragmenter.scala 109:20]
      end else begin
        r_addr_1 <= inc_addr_1; // @[Fragmenter.scala 107:35]
      end
    end
    r_len_1 <= _GEN_9[7:0];
    if (reset) begin // @[Fragmenter.scala 169:30]
      w_counter <= 9'h0; // @[Fragmenter.scala 169:30]
    end else begin
      w_counter <= _w_counter_T_2; // @[Fragmenter.scala 173:17]
    end
    if (reset) begin // @[Fragmenter.scala 155:35]
      wbeats_latched <= 1'h0; // @[Fragmenter.scala 155:35]
    end else if (_T_7) begin // @[Fragmenter.scala 159:26]
      wbeats_latched <= 1'h0; // @[Fragmenter.scala 159:43]
    end else begin
      wbeats_latched <= _GEN_10;
    end
    if (reset) begin // @[Fragmenter.scala 197:26]
      error_0 <= 2'h0; // @[Fragmenter.scala 197:26]
    end else if (_T_22[0] & _T_26) begin // @[Fragmenter.scala 200:34]
      if (auto_out_b_bits_echo_real_last) begin // @[Fragmenter.scala 200:46]
        error_0 <= 2'h0;
      end else begin
        error_0 <= _error_0_T;
      end
    end
    if (reset) begin // @[Fragmenter.scala 197:26]
      error_1 <= 2'h0; // @[Fragmenter.scala 197:26]
    end else if (_T_22[1] & _T_26) begin // @[Fragmenter.scala 200:34]
      if (auto_out_b_bits_echo_real_last) begin // @[Fragmenter.scala 200:46]
        error_1 <= 2'h0;
      end else begin
        error_1 <= _error_1_T;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~_w_counter_T | w_todo != 9'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Fragmenter.scala:174 assert (!out.w.fire || w_todo =/= 0.U) // underflow impossible\n"
            ); // @[Fragmenter.scala 174:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~_w_counter_T | w_todo != 9'h0) & ~reset) begin
          $fatal; // @[Fragmenter.scala 174:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & ~(~x1_w_valid | ~in_w_bits_last | w_last)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Fragmenter.scala:183 assert (!out.w.valid || !in_w.bits.last || w_last)\n"); // @[Fragmenter.scala 183:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~x1_w_valid | ~in_w_bits_last | w_last) & _T_13) begin
          $fatal; // @[Fragmenter.scala 183:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module AXI4IdIndexer_1(
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [15:0] auto_in_aw_bits_id,
  input  [15:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [1:0]  auto_in_aw_bits_burst,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [15:0] auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [15:0] auto_in_ar_bits_id,
  input  [15:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [1:0]  auto_in_ar_bits_burst,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [15:0] auto_in_r_bits_id,
  output [31:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output        auto_out_aw_bits_id,
  output [15:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  output [1:0]  auto_out_aw_bits_burst,
  output [14:0] auto_out_aw_bits_echo_extra_id,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [31:0] auto_out_w_bits_data,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input         auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input  [14:0] auto_out_b_bits_echo_extra_id,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output        auto_out_ar_bits_id,
  output [15:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output [1:0]  auto_out_ar_bits_burst,
  output [14:0] auto_out_ar_bits_echo_extra_id,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input         auto_out_r_bits_id,
  input  [31:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input  [14:0] auto_out_r_bits_echo_extra_id,
  input         auto_out_r_bits_last
);
  assign auto_in_aw_ready = auto_out_aw_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_w_ready = auto_out_w_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_b_valid = auto_out_b_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_b_bits_id = {auto_out_b_bits_echo_extra_id,auto_out_b_bits_id}; // @[Cat.scala 33:92]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_ar_ready = auto_out_ar_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_valid = auto_out_r_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_bits_id = {auto_out_r_bits_echo_extra_id,auto_out_r_bits_id}; // @[Cat.scala 33:92]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_r_bits_last = auto_out_r_bits_last; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_out_aw_valid = auto_in_aw_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id[0]; // @[Nodes.scala 1212:84 BundleMap.scala 247:19]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_len = auto_in_aw_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_size = auto_in_aw_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_burst = auto_in_aw_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_aw_bits_echo_extra_id = auto_in_aw_bits_id[15:1]; // @[IdIndexer.scala 74:56]
  assign auto_out_w_valid = auto_in_w_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_b_ready = auto_in_b_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_valid = auto_in_ar_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id[0]; // @[Nodes.scala 1212:84 BundleMap.scala 247:19]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_len = auto_in_ar_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_burst = auto_in_ar_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_ar_bits_echo_extra_id = auto_in_ar_bits_id[15:1]; // @[IdIndexer.scala 73:56]
  assign auto_out_r_ready = auto_in_r_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
endmodule
module Queue_180(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits
);
  reg [31:0] ram [0:15]; // @[Decoupled.scala 273:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [3:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [31:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [31:0] ram_MPORT_data; // @[Decoupled.scala 273:95]
  wire [3:0] ram_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 273:95]
  reg [3:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [3:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire [3:0] _value_T_1 = enq_ptr_value + 4'h1; // @[Counter.scala 77:24]
  wire [3:0] _value_T_3 = deq_ptr_value + 4'h1; // @[Counter.scala 77:24]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 4'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 4'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
endmodule
module Queue_181(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits
);
  reg [31:0] ram [0:15]; // @[Decoupled.scala 273:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [3:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [31:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [31:0] ram_MPORT_data; // @[Decoupled.scala 273:95]
  wire [3:0] ram_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 273:95]
  reg [3:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [3:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire [3:0] _value_T_1 = enq_ptr_value + 4'h1; // @[Counter.scala 77:24]
  wire [3:0] _value_T_3 = deq_ptr_value + 4'h1; // @[Counter.scala 77:24]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 4'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 4'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
endmodule
module AXILWidget(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [15:0] auto_in_aw_bits_id,
  input  [15:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [1:0]  auto_in_aw_bits_burst,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [15:0] auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [15:0] auto_in_ar_bits_id,
  input  [15:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [1:0]  auto_in_ar_bits_burst,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [15:0] auto_in_r_bits_id,
  output [31:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         io_cmds_ready,
  output        io_cmds_valid,
  output [31:0] io_cmds_bits,
  output        io_resp_ready,
  input         io_resp_valid,
  input  [31:0] io_resp_bits
);
  wire  crFile_clock; // @[AXILWidget.scala 13:35]
  wire  crFile_reset; // @[AXILWidget.scala 13:35]
  wire  crFile_auto_in_a_ready; // @[AXILWidget.scala 13:35]
  wire  crFile_auto_in_a_valid; // @[AXILWidget.scala 13:35]
  wire [2:0] crFile_auto_in_a_bits_opcode; // @[AXILWidget.scala 13:35]
  wire [3:0] crFile_auto_in_a_bits_source; // @[AXILWidget.scala 13:35]
  wire [15:0] crFile_auto_in_a_bits_address; // @[AXILWidget.scala 13:35]
  wire [31:0] crFile_auto_in_a_bits_data; // @[AXILWidget.scala 13:35]
  wire  crFile_auto_in_d_ready; // @[AXILWidget.scala 13:35]
  wire  crFile_auto_in_d_valid; // @[AXILWidget.scala 13:35]
  wire [2:0] crFile_auto_in_d_bits_opcode; // @[AXILWidget.scala 13:35]
  wire [3:0] crFile_auto_in_d_bits_source; // @[AXILWidget.scala 13:35]
  wire [31:0] crFile_auto_in_d_bits_data; // @[AXILWidget.scala 13:35]
  wire  crFile_io_mcr_read_0_ready; // @[AXILWidget.scala 13:35]
  wire [31:0] crFile_io_mcr_read_0_bits; // @[AXILWidget.scala 13:35]
  wire  crFile_io_mcr_read_1_ready; // @[AXILWidget.scala 13:35]
  wire [31:0] crFile_io_mcr_read_1_bits; // @[AXILWidget.scala 13:35]
  wire  crFile_io_mcr_read_2_ready; // @[AXILWidget.scala 13:35]
  wire [31:0] crFile_io_mcr_read_2_bits; // @[AXILWidget.scala 13:35]
  wire  crFile_io_mcr_read_3_ready; // @[AXILWidget.scala 13:35]
  wire [31:0] crFile_io_mcr_read_3_bits; // @[AXILWidget.scala 13:35]
  wire  crFile_io_mcr_read_4_ready; // @[AXILWidget.scala 13:35]
  wire [31:0] crFile_io_mcr_read_4_bits; // @[AXILWidget.scala 13:35]
  wire  crFile_io_mcr_read_5_ready; // @[AXILWidget.scala 13:35]
  wire [31:0] crFile_io_mcr_read_5_bits; // @[AXILWidget.scala 13:35]
  wire  crFile_io_mcr_read_6_ready; // @[AXILWidget.scala 13:35]
  wire [31:0] crFile_io_mcr_read_6_bits; // @[AXILWidget.scala 13:35]
  wire  crFile_io_mcr_read_7_ready; // @[AXILWidget.scala 13:35]
  wire  crFile_io_mcr_write_0_valid; // @[AXILWidget.scala 13:35]
  wire [31:0] crFile_io_mcr_write_0_bits; // @[AXILWidget.scala 13:35]
  wire  crFile_io_mcr_write_1_valid; // @[AXILWidget.scala 13:35]
  wire [31:0] crFile_io_mcr_write_1_bits; // @[AXILWidget.scala 13:35]
  wire  crFile_io_mcr_write_2_valid; // @[AXILWidget.scala 13:35]
  wire [31:0] crFile_io_mcr_write_2_bits; // @[AXILWidget.scala 13:35]
  wire  crFile_io_mcr_write_3_valid; // @[AXILWidget.scala 13:35]
  wire [31:0] crFile_io_mcr_write_3_bits; // @[AXILWidget.scala 13:35]
  wire  crFile_io_mcr_write_4_valid; // @[AXILWidget.scala 13:35]
  wire [31:0] crFile_io_mcr_write_4_bits; // @[AXILWidget.scala 13:35]
  wire  crFile_io_mcr_write_5_valid; // @[AXILWidget.scala 13:35]
  wire [31:0] crFile_io_mcr_write_5_bits; // @[AXILWidget.scala 13:35]
  wire  crFile_io_mcr_write_6_valid; // @[AXILWidget.scala 13:35]
  wire [31:0] crFile_io_mcr_write_6_bits; // @[AXILWidget.scala 13:35]
  wire  axi42tl_clock; // @[ToTL.scala 227:29]
  wire  axi42tl_reset; // @[ToTL.scala 227:29]
  wire  axi42tl_auto_in_aw_ready; // @[ToTL.scala 227:29]
  wire  axi42tl_auto_in_aw_valid; // @[ToTL.scala 227:29]
  wire  axi42tl_auto_in_aw_bits_id; // @[ToTL.scala 227:29]
  wire [15:0] axi42tl_auto_in_aw_bits_addr; // @[ToTL.scala 227:29]
  wire [2:0] axi42tl_auto_in_aw_bits_size; // @[ToTL.scala 227:29]
  wire  axi42tl_auto_in_w_ready; // @[ToTL.scala 227:29]
  wire  axi42tl_auto_in_w_valid; // @[ToTL.scala 227:29]
  wire [31:0] axi42tl_auto_in_w_bits_data; // @[ToTL.scala 227:29]
  wire  axi42tl_auto_in_w_bits_last; // @[ToTL.scala 227:29]
  wire  axi42tl_auto_in_b_ready; // @[ToTL.scala 227:29]
  wire  axi42tl_auto_in_b_valid; // @[ToTL.scala 227:29]
  wire  axi42tl_auto_in_b_bits_id; // @[ToTL.scala 227:29]
  wire [1:0] axi42tl_auto_in_b_bits_resp; // @[ToTL.scala 227:29]
  wire  axi42tl_auto_in_ar_ready; // @[ToTL.scala 227:29]
  wire  axi42tl_auto_in_ar_valid; // @[ToTL.scala 227:29]
  wire  axi42tl_auto_in_ar_bits_id; // @[ToTL.scala 227:29]
  wire [15:0] axi42tl_auto_in_ar_bits_addr; // @[ToTL.scala 227:29]
  wire [2:0] axi42tl_auto_in_ar_bits_size; // @[ToTL.scala 227:29]
  wire  axi42tl_auto_in_r_ready; // @[ToTL.scala 227:29]
  wire  axi42tl_auto_in_r_valid; // @[ToTL.scala 227:29]
  wire  axi42tl_auto_in_r_bits_id; // @[ToTL.scala 227:29]
  wire [31:0] axi42tl_auto_in_r_bits_data; // @[ToTL.scala 227:29]
  wire [1:0] axi42tl_auto_in_r_bits_resp; // @[ToTL.scala 227:29]
  wire  axi42tl_auto_in_r_bits_last; // @[ToTL.scala 227:29]
  wire  axi42tl_auto_out_a_ready; // @[ToTL.scala 227:29]
  wire  axi42tl_auto_out_a_valid; // @[ToTL.scala 227:29]
  wire [2:0] axi42tl_auto_out_a_bits_opcode; // @[ToTL.scala 227:29]
  wire [3:0] axi42tl_auto_out_a_bits_source; // @[ToTL.scala 227:29]
  wire [15:0] axi42tl_auto_out_a_bits_address; // @[ToTL.scala 227:29]
  wire [31:0] axi42tl_auto_out_a_bits_data; // @[ToTL.scala 227:29]
  wire  axi42tl_auto_out_d_ready; // @[ToTL.scala 227:29]
  wire  axi42tl_auto_out_d_valid; // @[ToTL.scala 227:29]
  wire [2:0] axi42tl_auto_out_d_bits_opcode; // @[ToTL.scala 227:29]
  wire [3:0] axi42tl_auto_out_d_bits_source; // @[ToTL.scala 227:29]
  wire [31:0] axi42tl_auto_out_d_bits_data; // @[ToTL.scala 227:29]
  wire  axi4yank_clock; // @[UserYanker.scala 108:30]
  wire  axi4yank_reset; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_aw_ready; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_aw_valid; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_aw_bits_id; // @[UserYanker.scala 108:30]
  wire [15:0] axi4yank_auto_in_aw_bits_addr; // @[UserYanker.scala 108:30]
  wire [2:0] axi4yank_auto_in_aw_bits_size; // @[UserYanker.scala 108:30]
  wire [14:0] axi4yank_auto_in_aw_bits_echo_extra_id; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_aw_bits_echo_real_last; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_w_ready; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_w_valid; // @[UserYanker.scala 108:30]
  wire [31:0] axi4yank_auto_in_w_bits_data; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_w_bits_last; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_b_ready; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_b_valid; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_b_bits_id; // @[UserYanker.scala 108:30]
  wire [1:0] axi4yank_auto_in_b_bits_resp; // @[UserYanker.scala 108:30]
  wire [14:0] axi4yank_auto_in_b_bits_echo_extra_id; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_b_bits_echo_real_last; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_ar_ready; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_ar_valid; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_ar_bits_id; // @[UserYanker.scala 108:30]
  wire [15:0] axi4yank_auto_in_ar_bits_addr; // @[UserYanker.scala 108:30]
  wire [2:0] axi4yank_auto_in_ar_bits_size; // @[UserYanker.scala 108:30]
  wire [14:0] axi4yank_auto_in_ar_bits_echo_extra_id; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_ar_bits_echo_real_last; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_r_ready; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_r_valid; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_r_bits_id; // @[UserYanker.scala 108:30]
  wire [31:0] axi4yank_auto_in_r_bits_data; // @[UserYanker.scala 108:30]
  wire [1:0] axi4yank_auto_in_r_bits_resp; // @[UserYanker.scala 108:30]
  wire [14:0] axi4yank_auto_in_r_bits_echo_extra_id; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_r_bits_echo_real_last; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_r_bits_last; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_aw_ready; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_aw_valid; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_aw_bits_id; // @[UserYanker.scala 108:30]
  wire [15:0] axi4yank_auto_out_aw_bits_addr; // @[UserYanker.scala 108:30]
  wire [2:0] axi4yank_auto_out_aw_bits_size; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_w_ready; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_w_valid; // @[UserYanker.scala 108:30]
  wire [31:0] axi4yank_auto_out_w_bits_data; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_w_bits_last; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_b_ready; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_b_valid; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_b_bits_id; // @[UserYanker.scala 108:30]
  wire [1:0] axi4yank_auto_out_b_bits_resp; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_ar_ready; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_ar_valid; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_ar_bits_id; // @[UserYanker.scala 108:30]
  wire [15:0] axi4yank_auto_out_ar_bits_addr; // @[UserYanker.scala 108:30]
  wire [2:0] axi4yank_auto_out_ar_bits_size; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_r_ready; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_r_valid; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_r_bits_id; // @[UserYanker.scala 108:30]
  wire [31:0] axi4yank_auto_out_r_bits_data; // @[UserYanker.scala 108:30]
  wire [1:0] axi4yank_auto_out_r_bits_resp; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_r_bits_last; // @[UserYanker.scala 108:30]
  wire  axi4frag_clock; // @[Fragmenter.scala 210:30]
  wire  axi4frag_reset; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_in_aw_ready; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_in_aw_valid; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_in_aw_bits_id; // @[Fragmenter.scala 210:30]
  wire [15:0] axi4frag_auto_in_aw_bits_addr; // @[Fragmenter.scala 210:30]
  wire [7:0] axi4frag_auto_in_aw_bits_len; // @[Fragmenter.scala 210:30]
  wire [2:0] axi4frag_auto_in_aw_bits_size; // @[Fragmenter.scala 210:30]
  wire [1:0] axi4frag_auto_in_aw_bits_burst; // @[Fragmenter.scala 210:30]
  wire [14:0] axi4frag_auto_in_aw_bits_echo_extra_id; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_in_w_ready; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_in_w_valid; // @[Fragmenter.scala 210:30]
  wire [31:0] axi4frag_auto_in_w_bits_data; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_in_w_bits_last; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_in_b_ready; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_in_b_valid; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_in_b_bits_id; // @[Fragmenter.scala 210:30]
  wire [1:0] axi4frag_auto_in_b_bits_resp; // @[Fragmenter.scala 210:30]
  wire [14:0] axi4frag_auto_in_b_bits_echo_extra_id; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_in_ar_ready; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_in_ar_valid; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_in_ar_bits_id; // @[Fragmenter.scala 210:30]
  wire [15:0] axi4frag_auto_in_ar_bits_addr; // @[Fragmenter.scala 210:30]
  wire [7:0] axi4frag_auto_in_ar_bits_len; // @[Fragmenter.scala 210:30]
  wire [2:0] axi4frag_auto_in_ar_bits_size; // @[Fragmenter.scala 210:30]
  wire [1:0] axi4frag_auto_in_ar_bits_burst; // @[Fragmenter.scala 210:30]
  wire [14:0] axi4frag_auto_in_ar_bits_echo_extra_id; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_in_r_ready; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_in_r_valid; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_in_r_bits_id; // @[Fragmenter.scala 210:30]
  wire [31:0] axi4frag_auto_in_r_bits_data; // @[Fragmenter.scala 210:30]
  wire [1:0] axi4frag_auto_in_r_bits_resp; // @[Fragmenter.scala 210:30]
  wire [14:0] axi4frag_auto_in_r_bits_echo_extra_id; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_in_r_bits_last; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_out_aw_ready; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_out_aw_valid; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_out_aw_bits_id; // @[Fragmenter.scala 210:30]
  wire [15:0] axi4frag_auto_out_aw_bits_addr; // @[Fragmenter.scala 210:30]
  wire [2:0] axi4frag_auto_out_aw_bits_size; // @[Fragmenter.scala 210:30]
  wire [14:0] axi4frag_auto_out_aw_bits_echo_extra_id; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_out_aw_bits_echo_real_last; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_out_w_ready; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_out_w_valid; // @[Fragmenter.scala 210:30]
  wire [31:0] axi4frag_auto_out_w_bits_data; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_out_w_bits_last; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_out_b_ready; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_out_b_valid; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_out_b_bits_id; // @[Fragmenter.scala 210:30]
  wire [1:0] axi4frag_auto_out_b_bits_resp; // @[Fragmenter.scala 210:30]
  wire [14:0] axi4frag_auto_out_b_bits_echo_extra_id; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_out_b_bits_echo_real_last; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_out_ar_ready; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_out_ar_valid; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_out_ar_bits_id; // @[Fragmenter.scala 210:30]
  wire [15:0] axi4frag_auto_out_ar_bits_addr; // @[Fragmenter.scala 210:30]
  wire [2:0] axi4frag_auto_out_ar_bits_size; // @[Fragmenter.scala 210:30]
  wire [14:0] axi4frag_auto_out_ar_bits_echo_extra_id; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_out_ar_bits_echo_real_last; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_out_r_ready; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_out_r_valid; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_out_r_bits_id; // @[Fragmenter.scala 210:30]
  wire [31:0] axi4frag_auto_out_r_bits_data; // @[Fragmenter.scala 210:30]
  wire [1:0] axi4frag_auto_out_r_bits_resp; // @[Fragmenter.scala 210:30]
  wire [14:0] axi4frag_auto_out_r_bits_echo_extra_id; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_out_r_bits_echo_real_last; // @[Fragmenter.scala 210:30]
  wire  axi4frag_auto_out_r_bits_last; // @[Fragmenter.scala 210:30]
  wire  axi4index_auto_in_aw_ready; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_in_aw_valid; // @[IdIndexer.scala 94:31]
  wire [15:0] axi4index_auto_in_aw_bits_id; // @[IdIndexer.scala 94:31]
  wire [15:0] axi4index_auto_in_aw_bits_addr; // @[IdIndexer.scala 94:31]
  wire [7:0] axi4index_auto_in_aw_bits_len; // @[IdIndexer.scala 94:31]
  wire [2:0] axi4index_auto_in_aw_bits_size; // @[IdIndexer.scala 94:31]
  wire [1:0] axi4index_auto_in_aw_bits_burst; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_in_w_ready; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_in_w_valid; // @[IdIndexer.scala 94:31]
  wire [31:0] axi4index_auto_in_w_bits_data; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_in_w_bits_last; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_in_b_ready; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_in_b_valid; // @[IdIndexer.scala 94:31]
  wire [15:0] axi4index_auto_in_b_bits_id; // @[IdIndexer.scala 94:31]
  wire [1:0] axi4index_auto_in_b_bits_resp; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_in_ar_ready; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_in_ar_valid; // @[IdIndexer.scala 94:31]
  wire [15:0] axi4index_auto_in_ar_bits_id; // @[IdIndexer.scala 94:31]
  wire [15:0] axi4index_auto_in_ar_bits_addr; // @[IdIndexer.scala 94:31]
  wire [7:0] axi4index_auto_in_ar_bits_len; // @[IdIndexer.scala 94:31]
  wire [2:0] axi4index_auto_in_ar_bits_size; // @[IdIndexer.scala 94:31]
  wire [1:0] axi4index_auto_in_ar_bits_burst; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_in_r_ready; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_in_r_valid; // @[IdIndexer.scala 94:31]
  wire [15:0] axi4index_auto_in_r_bits_id; // @[IdIndexer.scala 94:31]
  wire [31:0] axi4index_auto_in_r_bits_data; // @[IdIndexer.scala 94:31]
  wire [1:0] axi4index_auto_in_r_bits_resp; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_in_r_bits_last; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_aw_ready; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_aw_valid; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_aw_bits_id; // @[IdIndexer.scala 94:31]
  wire [15:0] axi4index_auto_out_aw_bits_addr; // @[IdIndexer.scala 94:31]
  wire [7:0] axi4index_auto_out_aw_bits_len; // @[IdIndexer.scala 94:31]
  wire [2:0] axi4index_auto_out_aw_bits_size; // @[IdIndexer.scala 94:31]
  wire [1:0] axi4index_auto_out_aw_bits_burst; // @[IdIndexer.scala 94:31]
  wire [14:0] axi4index_auto_out_aw_bits_echo_extra_id; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_w_ready; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_w_valid; // @[IdIndexer.scala 94:31]
  wire [31:0] axi4index_auto_out_w_bits_data; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_w_bits_last; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_b_ready; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_b_valid; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_b_bits_id; // @[IdIndexer.scala 94:31]
  wire [1:0] axi4index_auto_out_b_bits_resp; // @[IdIndexer.scala 94:31]
  wire [14:0] axi4index_auto_out_b_bits_echo_extra_id; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_ar_ready; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_ar_valid; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_ar_bits_id; // @[IdIndexer.scala 94:31]
  wire [15:0] axi4index_auto_out_ar_bits_addr; // @[IdIndexer.scala 94:31]
  wire [7:0] axi4index_auto_out_ar_bits_len; // @[IdIndexer.scala 94:31]
  wire [2:0] axi4index_auto_out_ar_bits_size; // @[IdIndexer.scala 94:31]
  wire [1:0] axi4index_auto_out_ar_bits_burst; // @[IdIndexer.scala 94:31]
  wire [14:0] axi4index_auto_out_ar_bits_echo_extra_id; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_r_ready; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_r_valid; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_r_bits_id; // @[IdIndexer.scala 94:31]
  wire [31:0] axi4index_auto_out_r_bits_data; // @[IdIndexer.scala 94:31]
  wire [1:0] axi4index_auto_out_r_bits_resp; // @[IdIndexer.scala 94:31]
  wire [14:0] axi4index_auto_out_r_bits_echo_extra_id; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_r_bits_last; // @[IdIndexer.scala 94:31]
  wire  roccCmdFifo_clock; // @[AXILWidget.scala 25:27]
  wire  roccCmdFifo_reset; // @[AXILWidget.scala 25:27]
  wire  roccCmdFifo_io_enq_ready; // @[AXILWidget.scala 25:27]
  wire  roccCmdFifo_io_enq_valid; // @[AXILWidget.scala 25:27]
  wire [31:0] roccCmdFifo_io_enq_bits; // @[AXILWidget.scala 25:27]
  wire  roccCmdFifo_io_deq_ready; // @[AXILWidget.scala 25:27]
  wire  roccCmdFifo_io_deq_valid; // @[AXILWidget.scala 25:27]
  wire [31:0] roccCmdFifo_io_deq_bits; // @[AXILWidget.scala 25:27]
  wire  roccRespFifo_clock; // @[AXILWidget.scala 26:28]
  wire  roccRespFifo_reset; // @[AXILWidget.scala 26:28]
  wire  roccRespFifo_io_enq_ready; // @[AXILWidget.scala 26:28]
  wire  roccRespFifo_io_enq_valid; // @[AXILWidget.scala 26:28]
  wire [31:0] roccRespFifo_io_enq_bits; // @[AXILWidget.scala 26:28]
  wire  roccRespFifo_io_deq_ready; // @[AXILWidget.scala 26:28]
  wire  roccRespFifo_io_deq_valid; // @[AXILWidget.scala 26:28]
  wire [31:0] roccRespFifo_io_deq_bits; // @[AXILWidget.scala 26:28]
  reg [31:0] resp_bits; // @[Widgets.scala 93:23]
  reg  resp_valid; // @[Widgets.scala 93:23]
  reg  resp_ready; // @[Widgets.scala 94:33]
  wire  _GEN_0 = resp_ready ? 1'h0 : resp_ready; // @[Widgets.scala 149:16 150:12 94:33]
  reg [31:0] cmd_bits; // @[Widgets.scala 93:23]
  reg  cmd_valid; // @[Widgets.scala 94:33]
  wire  _GEN_1 = cmd_valid ? 1'h0 : cmd_valid; // @[Widgets.scala 149:16 150:12 94:33]
  reg  cmd_ready; // @[Widgets.scala 93:23]
  reg [31:0] AXIL_DEBUG; // @[Widgets.scala 93:23]
  wire [31:0] _GEN_3 = crFile_io_mcr_write_1_valid ? crFile_io_mcr_write_1_bits : {{31'd0}, roccRespFifo_io_deq_valid}; // @[MCR.scala 83:31 84:18 Widgets.scala 96:44]
  wire [31:0] _GEN_4 = crFile_io_mcr_write_2_valid ? crFile_io_mcr_write_2_bits : {{31'd0}, _GEN_0}; // @[MCR.scala 83:31 84:18]
  wire [31:0] _GEN_6 = crFile_io_mcr_write_4_valid ? crFile_io_mcr_write_4_bits : {{31'd0}, _GEN_1}; // @[MCR.scala 83:31 84:18]
  wire [31:0] _GEN_7 = crFile_io_mcr_write_5_valid ? crFile_io_mcr_write_5_bits : {{31'd0}, roccCmdFifo_io_enq_ready}; // @[MCR.scala 83:31 84:18 Widgets.scala 96:44]
  wire [31:0] _GEN_9 = reset ? 32'h0 : _GEN_4; // @[Widgets.scala 94:{33,33}]
  wire [31:0] _GEN_10 = reset ? 32'h0 : _GEN_6; // @[Widgets.scala 94:{33,33}]
  MCRFileTL crFile ( // @[AXILWidget.scala 13:35]
    .clock(crFile_clock),
    .reset(crFile_reset),
    .auto_in_a_ready(crFile_auto_in_a_ready),
    .auto_in_a_valid(crFile_auto_in_a_valid),
    .auto_in_a_bits_opcode(crFile_auto_in_a_bits_opcode),
    .auto_in_a_bits_source(crFile_auto_in_a_bits_source),
    .auto_in_a_bits_address(crFile_auto_in_a_bits_address),
    .auto_in_a_bits_data(crFile_auto_in_a_bits_data),
    .auto_in_d_ready(crFile_auto_in_d_ready),
    .auto_in_d_valid(crFile_auto_in_d_valid),
    .auto_in_d_bits_opcode(crFile_auto_in_d_bits_opcode),
    .auto_in_d_bits_source(crFile_auto_in_d_bits_source),
    .auto_in_d_bits_data(crFile_auto_in_d_bits_data),
    .io_mcr_read_0_ready(crFile_io_mcr_read_0_ready),
    .io_mcr_read_0_bits(crFile_io_mcr_read_0_bits),
    .io_mcr_read_1_ready(crFile_io_mcr_read_1_ready),
    .io_mcr_read_1_bits(crFile_io_mcr_read_1_bits),
    .io_mcr_read_2_ready(crFile_io_mcr_read_2_ready),
    .io_mcr_read_2_bits(crFile_io_mcr_read_2_bits),
    .io_mcr_read_3_ready(crFile_io_mcr_read_3_ready),
    .io_mcr_read_3_bits(crFile_io_mcr_read_3_bits),
    .io_mcr_read_4_ready(crFile_io_mcr_read_4_ready),
    .io_mcr_read_4_bits(crFile_io_mcr_read_4_bits),
    .io_mcr_read_5_ready(crFile_io_mcr_read_5_ready),
    .io_mcr_read_5_bits(crFile_io_mcr_read_5_bits),
    .io_mcr_read_6_ready(crFile_io_mcr_read_6_ready),
    .io_mcr_read_6_bits(crFile_io_mcr_read_6_bits),
    .io_mcr_read_7_ready(crFile_io_mcr_read_7_ready),
    .io_mcr_write_0_valid(crFile_io_mcr_write_0_valid),
    .io_mcr_write_0_bits(crFile_io_mcr_write_0_bits),
    .io_mcr_write_1_valid(crFile_io_mcr_write_1_valid),
    .io_mcr_write_1_bits(crFile_io_mcr_write_1_bits),
    .io_mcr_write_2_valid(crFile_io_mcr_write_2_valid),
    .io_mcr_write_2_bits(crFile_io_mcr_write_2_bits),
    .io_mcr_write_3_valid(crFile_io_mcr_write_3_valid),
    .io_mcr_write_3_bits(crFile_io_mcr_write_3_bits),
    .io_mcr_write_4_valid(crFile_io_mcr_write_4_valid),
    .io_mcr_write_4_bits(crFile_io_mcr_write_4_bits),
    .io_mcr_write_5_valid(crFile_io_mcr_write_5_valid),
    .io_mcr_write_5_bits(crFile_io_mcr_write_5_bits),
    .io_mcr_write_6_valid(crFile_io_mcr_write_6_valid),
    .io_mcr_write_6_bits(crFile_io_mcr_write_6_bits)
  );
  AXI4ToTL axi42tl ( // @[ToTL.scala 227:29]
    .clock(axi42tl_clock),
    .reset(axi42tl_reset),
    .auto_in_aw_ready(axi42tl_auto_in_aw_ready),
    .auto_in_aw_valid(axi42tl_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi42tl_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi42tl_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi42tl_auto_in_aw_bits_size),
    .auto_in_w_ready(axi42tl_auto_in_w_ready),
    .auto_in_w_valid(axi42tl_auto_in_w_valid),
    .auto_in_w_bits_data(axi42tl_auto_in_w_bits_data),
    .auto_in_w_bits_last(axi42tl_auto_in_w_bits_last),
    .auto_in_b_ready(axi42tl_auto_in_b_ready),
    .auto_in_b_valid(axi42tl_auto_in_b_valid),
    .auto_in_b_bits_id(axi42tl_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi42tl_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi42tl_auto_in_ar_ready),
    .auto_in_ar_valid(axi42tl_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi42tl_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi42tl_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi42tl_auto_in_ar_bits_size),
    .auto_in_r_ready(axi42tl_auto_in_r_ready),
    .auto_in_r_valid(axi42tl_auto_in_r_valid),
    .auto_in_r_bits_id(axi42tl_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi42tl_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi42tl_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi42tl_auto_in_r_bits_last),
    .auto_out_a_ready(axi42tl_auto_out_a_ready),
    .auto_out_a_valid(axi42tl_auto_out_a_valid),
    .auto_out_a_bits_opcode(axi42tl_auto_out_a_bits_opcode),
    .auto_out_a_bits_source(axi42tl_auto_out_a_bits_source),
    .auto_out_a_bits_address(axi42tl_auto_out_a_bits_address),
    .auto_out_a_bits_data(axi42tl_auto_out_a_bits_data),
    .auto_out_d_ready(axi42tl_auto_out_d_ready),
    .auto_out_d_valid(axi42tl_auto_out_d_valid),
    .auto_out_d_bits_opcode(axi42tl_auto_out_d_bits_opcode),
    .auto_out_d_bits_source(axi42tl_auto_out_d_bits_source),
    .auto_out_d_bits_data(axi42tl_auto_out_d_bits_data)
  );
  AXI4UserYanker_1 axi4yank ( // @[UserYanker.scala 108:30]
    .clock(axi4yank_clock),
    .reset(axi4yank_reset),
    .auto_in_aw_ready(axi4yank_auto_in_aw_ready),
    .auto_in_aw_valid(axi4yank_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4yank_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4yank_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4yank_auto_in_aw_bits_size),
    .auto_in_aw_bits_echo_extra_id(axi4yank_auto_in_aw_bits_echo_extra_id),
    .auto_in_aw_bits_echo_real_last(axi4yank_auto_in_aw_bits_echo_real_last),
    .auto_in_w_ready(axi4yank_auto_in_w_ready),
    .auto_in_w_valid(axi4yank_auto_in_w_valid),
    .auto_in_w_bits_data(axi4yank_auto_in_w_bits_data),
    .auto_in_w_bits_last(axi4yank_auto_in_w_bits_last),
    .auto_in_b_ready(axi4yank_auto_in_b_ready),
    .auto_in_b_valid(axi4yank_auto_in_b_valid),
    .auto_in_b_bits_id(axi4yank_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4yank_auto_in_b_bits_resp),
    .auto_in_b_bits_echo_extra_id(axi4yank_auto_in_b_bits_echo_extra_id),
    .auto_in_b_bits_echo_real_last(axi4yank_auto_in_b_bits_echo_real_last),
    .auto_in_ar_ready(axi4yank_auto_in_ar_ready),
    .auto_in_ar_valid(axi4yank_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4yank_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4yank_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4yank_auto_in_ar_bits_size),
    .auto_in_ar_bits_echo_extra_id(axi4yank_auto_in_ar_bits_echo_extra_id),
    .auto_in_ar_bits_echo_real_last(axi4yank_auto_in_ar_bits_echo_real_last),
    .auto_in_r_ready(axi4yank_auto_in_r_ready),
    .auto_in_r_valid(axi4yank_auto_in_r_valid),
    .auto_in_r_bits_id(axi4yank_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4yank_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4yank_auto_in_r_bits_resp),
    .auto_in_r_bits_echo_extra_id(axi4yank_auto_in_r_bits_echo_extra_id),
    .auto_in_r_bits_echo_real_last(axi4yank_auto_in_r_bits_echo_real_last),
    .auto_in_r_bits_last(axi4yank_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4yank_auto_out_aw_ready),
    .auto_out_aw_valid(axi4yank_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4yank_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4yank_auto_out_aw_bits_addr),
    .auto_out_aw_bits_size(axi4yank_auto_out_aw_bits_size),
    .auto_out_w_ready(axi4yank_auto_out_w_ready),
    .auto_out_w_valid(axi4yank_auto_out_w_valid),
    .auto_out_w_bits_data(axi4yank_auto_out_w_bits_data),
    .auto_out_w_bits_last(axi4yank_auto_out_w_bits_last),
    .auto_out_b_ready(axi4yank_auto_out_b_ready),
    .auto_out_b_valid(axi4yank_auto_out_b_valid),
    .auto_out_b_bits_id(axi4yank_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4yank_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4yank_auto_out_ar_ready),
    .auto_out_ar_valid(axi4yank_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4yank_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4yank_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4yank_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4yank_auto_out_r_ready),
    .auto_out_r_valid(axi4yank_auto_out_r_valid),
    .auto_out_r_bits_id(axi4yank_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4yank_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4yank_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4yank_auto_out_r_bits_last)
  );
  AXI4Fragmenter axi4frag ( // @[Fragmenter.scala 210:30]
    .clock(axi4frag_clock),
    .reset(axi4frag_reset),
    .auto_in_aw_ready(axi4frag_auto_in_aw_ready),
    .auto_in_aw_valid(axi4frag_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4frag_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4frag_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4frag_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4frag_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axi4frag_auto_in_aw_bits_burst),
    .auto_in_aw_bits_echo_extra_id(axi4frag_auto_in_aw_bits_echo_extra_id),
    .auto_in_w_ready(axi4frag_auto_in_w_ready),
    .auto_in_w_valid(axi4frag_auto_in_w_valid),
    .auto_in_w_bits_data(axi4frag_auto_in_w_bits_data),
    .auto_in_w_bits_last(axi4frag_auto_in_w_bits_last),
    .auto_in_b_ready(axi4frag_auto_in_b_ready),
    .auto_in_b_valid(axi4frag_auto_in_b_valid),
    .auto_in_b_bits_id(axi4frag_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4frag_auto_in_b_bits_resp),
    .auto_in_b_bits_echo_extra_id(axi4frag_auto_in_b_bits_echo_extra_id),
    .auto_in_ar_ready(axi4frag_auto_in_ar_ready),
    .auto_in_ar_valid(axi4frag_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4frag_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4frag_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4frag_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4frag_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axi4frag_auto_in_ar_bits_burst),
    .auto_in_ar_bits_echo_extra_id(axi4frag_auto_in_ar_bits_echo_extra_id),
    .auto_in_r_ready(axi4frag_auto_in_r_ready),
    .auto_in_r_valid(axi4frag_auto_in_r_valid),
    .auto_in_r_bits_id(axi4frag_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4frag_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4frag_auto_in_r_bits_resp),
    .auto_in_r_bits_echo_extra_id(axi4frag_auto_in_r_bits_echo_extra_id),
    .auto_in_r_bits_last(axi4frag_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4frag_auto_out_aw_ready),
    .auto_out_aw_valid(axi4frag_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4frag_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4frag_auto_out_aw_bits_addr),
    .auto_out_aw_bits_size(axi4frag_auto_out_aw_bits_size),
    .auto_out_aw_bits_echo_extra_id(axi4frag_auto_out_aw_bits_echo_extra_id),
    .auto_out_aw_bits_echo_real_last(axi4frag_auto_out_aw_bits_echo_real_last),
    .auto_out_w_ready(axi4frag_auto_out_w_ready),
    .auto_out_w_valid(axi4frag_auto_out_w_valid),
    .auto_out_w_bits_data(axi4frag_auto_out_w_bits_data),
    .auto_out_w_bits_last(axi4frag_auto_out_w_bits_last),
    .auto_out_b_ready(axi4frag_auto_out_b_ready),
    .auto_out_b_valid(axi4frag_auto_out_b_valid),
    .auto_out_b_bits_id(axi4frag_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4frag_auto_out_b_bits_resp),
    .auto_out_b_bits_echo_extra_id(axi4frag_auto_out_b_bits_echo_extra_id),
    .auto_out_b_bits_echo_real_last(axi4frag_auto_out_b_bits_echo_real_last),
    .auto_out_ar_ready(axi4frag_auto_out_ar_ready),
    .auto_out_ar_valid(axi4frag_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4frag_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4frag_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4frag_auto_out_ar_bits_size),
    .auto_out_ar_bits_echo_extra_id(axi4frag_auto_out_ar_bits_echo_extra_id),
    .auto_out_ar_bits_echo_real_last(axi4frag_auto_out_ar_bits_echo_real_last),
    .auto_out_r_ready(axi4frag_auto_out_r_ready),
    .auto_out_r_valid(axi4frag_auto_out_r_valid),
    .auto_out_r_bits_id(axi4frag_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4frag_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4frag_auto_out_r_bits_resp),
    .auto_out_r_bits_echo_extra_id(axi4frag_auto_out_r_bits_echo_extra_id),
    .auto_out_r_bits_echo_real_last(axi4frag_auto_out_r_bits_echo_real_last),
    .auto_out_r_bits_last(axi4frag_auto_out_r_bits_last)
  );
  AXI4IdIndexer_1 axi4index ( // @[IdIndexer.scala 94:31]
    .auto_in_aw_ready(axi4index_auto_in_aw_ready),
    .auto_in_aw_valid(axi4index_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4index_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4index_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4index_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4index_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axi4index_auto_in_aw_bits_burst),
    .auto_in_w_ready(axi4index_auto_in_w_ready),
    .auto_in_w_valid(axi4index_auto_in_w_valid),
    .auto_in_w_bits_data(axi4index_auto_in_w_bits_data),
    .auto_in_w_bits_last(axi4index_auto_in_w_bits_last),
    .auto_in_b_ready(axi4index_auto_in_b_ready),
    .auto_in_b_valid(axi4index_auto_in_b_valid),
    .auto_in_b_bits_id(axi4index_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4index_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4index_auto_in_ar_ready),
    .auto_in_ar_valid(axi4index_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4index_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4index_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4index_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4index_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axi4index_auto_in_ar_bits_burst),
    .auto_in_r_ready(axi4index_auto_in_r_ready),
    .auto_in_r_valid(axi4index_auto_in_r_valid),
    .auto_in_r_bits_id(axi4index_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4index_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4index_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4index_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4index_auto_out_aw_ready),
    .auto_out_aw_valid(axi4index_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4index_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4index_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4index_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4index_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(axi4index_auto_out_aw_bits_burst),
    .auto_out_aw_bits_echo_extra_id(axi4index_auto_out_aw_bits_echo_extra_id),
    .auto_out_w_ready(axi4index_auto_out_w_ready),
    .auto_out_w_valid(axi4index_auto_out_w_valid),
    .auto_out_w_bits_data(axi4index_auto_out_w_bits_data),
    .auto_out_w_bits_last(axi4index_auto_out_w_bits_last),
    .auto_out_b_ready(axi4index_auto_out_b_ready),
    .auto_out_b_valid(axi4index_auto_out_b_valid),
    .auto_out_b_bits_id(axi4index_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4index_auto_out_b_bits_resp),
    .auto_out_b_bits_echo_extra_id(axi4index_auto_out_b_bits_echo_extra_id),
    .auto_out_ar_ready(axi4index_auto_out_ar_ready),
    .auto_out_ar_valid(axi4index_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4index_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4index_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4index_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4index_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(axi4index_auto_out_ar_bits_burst),
    .auto_out_ar_bits_echo_extra_id(axi4index_auto_out_ar_bits_echo_extra_id),
    .auto_out_r_ready(axi4index_auto_out_r_ready),
    .auto_out_r_valid(axi4index_auto_out_r_valid),
    .auto_out_r_bits_id(axi4index_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4index_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4index_auto_out_r_bits_resp),
    .auto_out_r_bits_echo_extra_id(axi4index_auto_out_r_bits_echo_extra_id),
    .auto_out_r_bits_last(axi4index_auto_out_r_bits_last)
  );
  Queue_180 roccCmdFifo ( // @[AXILWidget.scala 25:27]
    .clock(roccCmdFifo_clock),
    .reset(roccCmdFifo_reset),
    .io_enq_ready(roccCmdFifo_io_enq_ready),
    .io_enq_valid(roccCmdFifo_io_enq_valid),
    .io_enq_bits(roccCmdFifo_io_enq_bits),
    .io_deq_ready(roccCmdFifo_io_deq_ready),
    .io_deq_valid(roccCmdFifo_io_deq_valid),
    .io_deq_bits(roccCmdFifo_io_deq_bits)
  );
  Queue_181 roccRespFifo ( // @[AXILWidget.scala 26:28]
    .clock(roccRespFifo_clock),
    .reset(roccRespFifo_reset),
    .io_enq_ready(roccRespFifo_io_enq_ready),
    .io_enq_valid(roccRespFifo_io_enq_valid),
    .io_enq_bits(roccRespFifo_io_enq_bits),
    .io_deq_ready(roccRespFifo_io_deq_ready),
    .io_deq_valid(roccRespFifo_io_deq_valid),
    .io_deq_bits(roccRespFifo_io_deq_bits)
  );
  assign auto_in_aw_ready = axi4index_auto_in_aw_ready; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign auto_in_w_ready = axi4index_auto_in_w_ready; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign auto_in_b_valid = axi4index_auto_in_b_valid; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign auto_in_b_bits_id = axi4index_auto_in_b_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign auto_in_b_bits_resp = axi4index_auto_in_b_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign auto_in_ar_ready = axi4index_auto_in_ar_ready; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign auto_in_r_valid = axi4index_auto_in_r_valid; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign auto_in_r_bits_id = axi4index_auto_in_r_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign auto_in_r_bits_data = axi4index_auto_in_r_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign auto_in_r_bits_resp = axi4index_auto_in_r_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign auto_in_r_bits_last = axi4index_auto_in_r_bits_last; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign io_cmds_valid = roccCmdFifo_io_deq_valid; // @[AXILWidget.scala 40:11]
  assign io_cmds_bits = roccCmdFifo_io_deq_bits; // @[AXILWidget.scala 40:11]
  assign io_resp_ready = roccRespFifo_io_enq_ready; // @[AXILWidget.scala 41:23]
  assign crFile_clock = clock;
  assign crFile_reset = reset;
  assign crFile_auto_in_a_valid = axi42tl_auto_out_a_valid; // @[LazyModule.scala 353:16]
  assign crFile_auto_in_a_bits_opcode = axi42tl_auto_out_a_bits_opcode; // @[LazyModule.scala 353:16]
  assign crFile_auto_in_a_bits_source = axi42tl_auto_out_a_bits_source; // @[LazyModule.scala 353:16]
  assign crFile_auto_in_a_bits_address = axi42tl_auto_out_a_bits_address; // @[LazyModule.scala 353:16]
  assign crFile_auto_in_a_bits_data = axi42tl_auto_out_a_bits_data; // @[LazyModule.scala 353:16]
  assign crFile_auto_in_d_ready = axi42tl_auto_out_d_ready; // @[LazyModule.scala 353:16]
  assign crFile_io_mcr_read_0_bits = resp_bits; // @[MCR.scala 91:23]
  assign crFile_io_mcr_read_1_bits = {{31'd0}, resp_valid}; // @[MCR.scala 91:23]
  assign crFile_io_mcr_read_2_bits = {{31'd0}, resp_ready}; // @[MCR.scala 91:23]
  assign crFile_io_mcr_read_3_bits = cmd_bits; // @[MCR.scala 91:23]
  assign crFile_io_mcr_read_4_bits = {{31'd0}, cmd_valid}; // @[MCR.scala 91:23]
  assign crFile_io_mcr_read_5_bits = {{31'd0}, cmd_ready}; // @[MCR.scala 91:23]
  assign crFile_io_mcr_read_6_bits = AXIL_DEBUG; // @[MCR.scala 91:23]
  assign axi42tl_clock = clock;
  assign axi42tl_reset = reset;
  assign axi42tl_auto_in_aw_valid = axi4yank_auto_out_aw_valid; // @[LazyModule.scala 353:16]
  assign axi42tl_auto_in_aw_bits_id = axi4yank_auto_out_aw_bits_id; // @[LazyModule.scala 353:16]
  assign axi42tl_auto_in_aw_bits_addr = axi4yank_auto_out_aw_bits_addr; // @[LazyModule.scala 353:16]
  assign axi42tl_auto_in_aw_bits_size = axi4yank_auto_out_aw_bits_size; // @[LazyModule.scala 353:16]
  assign axi42tl_auto_in_w_valid = axi4yank_auto_out_w_valid; // @[LazyModule.scala 353:16]
  assign axi42tl_auto_in_w_bits_data = axi4yank_auto_out_w_bits_data; // @[LazyModule.scala 353:16]
  assign axi42tl_auto_in_w_bits_last = axi4yank_auto_out_w_bits_last; // @[LazyModule.scala 353:16]
  assign axi42tl_auto_in_b_ready = axi4yank_auto_out_b_ready; // @[LazyModule.scala 353:16]
  assign axi42tl_auto_in_ar_valid = axi4yank_auto_out_ar_valid; // @[LazyModule.scala 353:16]
  assign axi42tl_auto_in_ar_bits_id = axi4yank_auto_out_ar_bits_id; // @[LazyModule.scala 353:16]
  assign axi42tl_auto_in_ar_bits_addr = axi4yank_auto_out_ar_bits_addr; // @[LazyModule.scala 353:16]
  assign axi42tl_auto_in_ar_bits_size = axi4yank_auto_out_ar_bits_size; // @[LazyModule.scala 353:16]
  assign axi42tl_auto_in_r_ready = axi4yank_auto_out_r_ready; // @[LazyModule.scala 353:16]
  assign axi42tl_auto_out_a_ready = crFile_auto_in_a_ready; // @[LazyModule.scala 353:16]
  assign axi42tl_auto_out_d_valid = crFile_auto_in_d_valid; // @[LazyModule.scala 353:16]
  assign axi42tl_auto_out_d_bits_opcode = crFile_auto_in_d_bits_opcode; // @[LazyModule.scala 353:16]
  assign axi42tl_auto_out_d_bits_source = crFile_auto_in_d_bits_source; // @[LazyModule.scala 353:16]
  assign axi42tl_auto_out_d_bits_data = crFile_auto_in_d_bits_data; // @[LazyModule.scala 353:16]
  assign axi4yank_clock = clock;
  assign axi4yank_reset = reset;
  assign axi4yank_auto_in_aw_valid = axi4frag_auto_out_aw_valid; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_aw_bits_id = axi4frag_auto_out_aw_bits_id; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_aw_bits_addr = axi4frag_auto_out_aw_bits_addr; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_aw_bits_size = axi4frag_auto_out_aw_bits_size; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_aw_bits_echo_extra_id = axi4frag_auto_out_aw_bits_echo_extra_id; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_aw_bits_echo_real_last = axi4frag_auto_out_aw_bits_echo_real_last; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_w_valid = axi4frag_auto_out_w_valid; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_w_bits_data = axi4frag_auto_out_w_bits_data; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_w_bits_last = axi4frag_auto_out_w_bits_last; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_b_ready = axi4frag_auto_out_b_ready; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_ar_valid = axi4frag_auto_out_ar_valid; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_ar_bits_id = axi4frag_auto_out_ar_bits_id; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_ar_bits_addr = axi4frag_auto_out_ar_bits_addr; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_ar_bits_size = axi4frag_auto_out_ar_bits_size; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_ar_bits_echo_extra_id = axi4frag_auto_out_ar_bits_echo_extra_id; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_ar_bits_echo_real_last = axi4frag_auto_out_ar_bits_echo_real_last; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_r_ready = axi4frag_auto_out_r_ready; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_out_aw_ready = axi42tl_auto_in_aw_ready; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_out_w_ready = axi42tl_auto_in_w_ready; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_out_b_valid = axi42tl_auto_in_b_valid; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_out_b_bits_id = axi42tl_auto_in_b_bits_id; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_out_b_bits_resp = axi42tl_auto_in_b_bits_resp; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_out_ar_ready = axi42tl_auto_in_ar_ready; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_out_r_valid = axi42tl_auto_in_r_valid; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_out_r_bits_id = axi42tl_auto_in_r_bits_id; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_out_r_bits_data = axi42tl_auto_in_r_bits_data; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_out_r_bits_resp = axi42tl_auto_in_r_bits_resp; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_out_r_bits_last = axi42tl_auto_in_r_bits_last; // @[LazyModule.scala 353:16]
  assign axi4frag_clock = clock;
  assign axi4frag_reset = reset;
  assign axi4frag_auto_in_aw_valid = axi4index_auto_out_aw_valid; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_in_aw_bits_id = axi4index_auto_out_aw_bits_id; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_in_aw_bits_addr = axi4index_auto_out_aw_bits_addr; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_in_aw_bits_len = axi4index_auto_out_aw_bits_len; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_in_aw_bits_size = axi4index_auto_out_aw_bits_size; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_in_aw_bits_burst = axi4index_auto_out_aw_bits_burst; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_in_aw_bits_echo_extra_id = axi4index_auto_out_aw_bits_echo_extra_id; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_in_w_valid = axi4index_auto_out_w_valid; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_in_w_bits_data = axi4index_auto_out_w_bits_data; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_in_w_bits_last = axi4index_auto_out_w_bits_last; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_in_b_ready = axi4index_auto_out_b_ready; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_in_ar_valid = axi4index_auto_out_ar_valid; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_in_ar_bits_id = axi4index_auto_out_ar_bits_id; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_in_ar_bits_addr = axi4index_auto_out_ar_bits_addr; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_in_ar_bits_len = axi4index_auto_out_ar_bits_len; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_in_ar_bits_size = axi4index_auto_out_ar_bits_size; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_in_ar_bits_burst = axi4index_auto_out_ar_bits_burst; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_in_ar_bits_echo_extra_id = axi4index_auto_out_ar_bits_echo_extra_id; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_in_r_ready = axi4index_auto_out_r_ready; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_out_aw_ready = axi4yank_auto_in_aw_ready; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_out_w_ready = axi4yank_auto_in_w_ready; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_out_b_valid = axi4yank_auto_in_b_valid; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_out_b_bits_id = axi4yank_auto_in_b_bits_id; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_out_b_bits_resp = axi4yank_auto_in_b_bits_resp; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_out_b_bits_echo_extra_id = axi4yank_auto_in_b_bits_echo_extra_id; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_out_b_bits_echo_real_last = axi4yank_auto_in_b_bits_echo_real_last; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_out_ar_ready = axi4yank_auto_in_ar_ready; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_out_r_valid = axi4yank_auto_in_r_valid; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_out_r_bits_id = axi4yank_auto_in_r_bits_id; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_out_r_bits_data = axi4yank_auto_in_r_bits_data; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_out_r_bits_resp = axi4yank_auto_in_r_bits_resp; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_out_r_bits_echo_extra_id = axi4yank_auto_in_r_bits_echo_extra_id; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_out_r_bits_echo_real_last = axi4yank_auto_in_r_bits_echo_real_last; // @[LazyModule.scala 353:16]
  assign axi4frag_auto_out_r_bits_last = axi4yank_auto_in_r_bits_last; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_aw_valid = auto_in_aw_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axi4index_auto_in_aw_bits_id = auto_in_aw_bits_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axi4index_auto_in_aw_bits_addr = auto_in_aw_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axi4index_auto_in_aw_bits_len = auto_in_aw_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axi4index_auto_in_aw_bits_size = auto_in_aw_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axi4index_auto_in_aw_bits_burst = auto_in_aw_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axi4index_auto_in_w_valid = auto_in_w_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axi4index_auto_in_w_bits_data = auto_in_w_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axi4index_auto_in_w_bits_last = auto_in_w_bits_last; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axi4index_auto_in_b_ready = auto_in_b_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axi4index_auto_in_ar_valid = auto_in_ar_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axi4index_auto_in_ar_bits_id = auto_in_ar_bits_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axi4index_auto_in_ar_bits_addr = auto_in_ar_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axi4index_auto_in_ar_bits_len = auto_in_ar_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axi4index_auto_in_ar_bits_size = auto_in_ar_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axi4index_auto_in_ar_bits_burst = auto_in_ar_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axi4index_auto_in_r_ready = auto_in_r_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axi4index_auto_out_aw_ready = axi4frag_auto_in_aw_ready; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_w_ready = axi4frag_auto_in_w_ready; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_b_valid = axi4frag_auto_in_b_valid; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_b_bits_id = axi4frag_auto_in_b_bits_id; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_b_bits_resp = axi4frag_auto_in_b_bits_resp; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_b_bits_echo_extra_id = axi4frag_auto_in_b_bits_echo_extra_id; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_ar_ready = axi4frag_auto_in_ar_ready; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_r_valid = axi4frag_auto_in_r_valid; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_r_bits_id = axi4frag_auto_in_r_bits_id; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_r_bits_data = axi4frag_auto_in_r_bits_data; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_r_bits_resp = axi4frag_auto_in_r_bits_resp; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_r_bits_echo_extra_id = axi4frag_auto_in_r_bits_echo_extra_id; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_r_bits_last = axi4frag_auto_in_r_bits_last; // @[LazyModule.scala 353:16]
  assign roccCmdFifo_clock = clock;
  assign roccCmdFifo_reset = reset;
  assign roccCmdFifo_io_enq_valid = cmd_valid; // @[Widgets.scala 96:28]
  assign roccCmdFifo_io_enq_bits = cmd_bits; // @[Widgets.scala 96:28]
  assign roccCmdFifo_io_deq_ready = io_cmds_ready; // @[AXILWidget.scala 40:11]
  assign roccRespFifo_clock = clock;
  assign roccRespFifo_reset = reset;
  assign roccRespFifo_io_enq_valid = io_resp_valid; // @[AXILWidget.scala 41:23]
  assign roccRespFifo_io_enq_bits = io_resp_bits; // @[AXILWidget.scala 41:23]
  assign roccRespFifo_io_deq_ready = resp_ready; // @[Widgets.scala 96:28]
  always @(posedge clock) begin
    if (crFile_io_mcr_write_0_valid) begin // @[MCR.scala 83:31]
      resp_bits <= crFile_io_mcr_write_0_bits; // @[MCR.scala 84:18]
    end else begin
      resp_bits <= roccRespFifo_io_deq_bits; // @[Widgets.scala 96:44]
    end
    resp_valid <= _GEN_3[0];
    resp_ready <= _GEN_9[0]; // @[Widgets.scala 94:{33,33}]
    if (crFile_io_mcr_write_3_valid) begin // @[MCR.scala 83:31]
      cmd_bits <= crFile_io_mcr_write_3_bits; // @[MCR.scala 84:18]
    end
    cmd_valid <= _GEN_10[0]; // @[Widgets.scala 94:{33,33}]
    cmd_ready <= _GEN_7[0];
    if (crFile_io_mcr_write_6_valid) begin // @[MCR.scala 83:31]
      AXIL_DEBUG <= crFile_io_mcr_write_6_bits; // @[MCR.scala 84:18]
    end else begin
      AXIL_DEBUG <= 32'hdeadcafe; // @[Widgets.scala 96:44]
    end
  end
endmodule
module AXILToRocc(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits,
  input         io_rocc_ready,
  output        io_rocc_valid,
  output [6:0]  io_rocc_bits_inst_funct,
  output [4:0]  io_rocc_bits_inst_rs2,
  output [4:0]  io_rocc_bits_inst_rs1,
  output [6:0]  io_rocc_bits_inst_opcode,
  output [63:0] io_rocc_bits_rs1,
  output [63:0] io_rocc_bits_rs2
);
  reg [3:0] counter; // @[AXILToRocc.scala 24:24]
  reg [31:0] bitsBuffer_0; // @[AXILToRocc.scala 25:23]
  reg [31:0] bitsBuffer_1; // @[AXILToRocc.scala 25:23]
  reg [31:0] bitsBuffer_2; // @[AXILToRocc.scala 25:23]
  reg [31:0] bitsBuffer_3; // @[AXILToRocc.scala 25:23]
  reg [31:0] bitsBuffer_4; // @[AXILToRocc.scala 25:23]
  wire  _T = io_in_ready & io_in_valid; // @[Decoupled.scala 51:35]
  wire [3:0] _counter_T_1 = counter + 4'h1; // @[AXILToRocc.scala 38:24]
  wire  _T_2 = io_rocc_ready & io_rocc_valid; // @[Decoupled.scala 51:35]
  assign io_in_ready = counter < 4'h5 & io_rocc_ready; // @[AXILToRocc.scala 34:39]
  assign io_rocc_valid = counter == 4'h5; // @[AXILToRocc.scala 35:29]
  assign io_rocc_bits_inst_funct = bitsBuffer_0[31:25]; // @[AXILToRocc.scala 29:38]
  assign io_rocc_bits_inst_rs2 = bitsBuffer_0[24:20]; // @[AXILToRocc.scala 29:38]
  assign io_rocc_bits_inst_rs1 = bitsBuffer_0[19:15]; // @[AXILToRocc.scala 29:38]
  assign io_rocc_bits_inst_opcode = bitsBuffer_0[6:0]; // @[AXILToRocc.scala 29:38]
  assign io_rocc_bits_rs1 = {bitsBuffer_1,bitsBuffer_2}; // @[Cat.scala 33:92]
  assign io_rocc_bits_rs2 = {bitsBuffer_3,bitsBuffer_4}; // @[Cat.scala 33:92]
  always @(posedge clock) begin
    if (reset) begin // @[AXILToRocc.scala 24:24]
      counter <= 4'h0; // @[AXILToRocc.scala 24:24]
    end else if (_T_2) begin // @[AXILToRocc.scala 41:22]
      counter <= 4'h0; // @[AXILToRocc.scala 42:13]
    end else if (_T) begin // @[AXILToRocc.scala 36:20]
      counter <= _counter_T_1; // @[AXILToRocc.scala 38:13]
    end
    if (_T) begin // @[AXILToRocc.scala 36:20]
      if (3'h0 == counter[2:0]) begin // @[AXILToRocc.scala 37:25]
        bitsBuffer_0 <= io_in_bits; // @[AXILToRocc.scala 37:25]
      end
    end
    if (_T) begin // @[AXILToRocc.scala 36:20]
      if (3'h1 == counter[2:0]) begin // @[AXILToRocc.scala 37:25]
        bitsBuffer_1 <= io_in_bits; // @[AXILToRocc.scala 37:25]
      end
    end
    if (_T) begin // @[AXILToRocc.scala 36:20]
      if (3'h2 == counter[2:0]) begin // @[AXILToRocc.scala 37:25]
        bitsBuffer_2 <= io_in_bits; // @[AXILToRocc.scala 37:25]
      end
    end
    if (_T) begin // @[AXILToRocc.scala 36:20]
      if (3'h3 == counter[2:0]) begin // @[AXILToRocc.scala 37:25]
        bitsBuffer_3 <= io_in_bits; // @[AXILToRocc.scala 37:25]
      end
    end
    if (_T) begin // @[AXILToRocc.scala 36:20]
      if (3'h4 == counter[2:0]) begin // @[AXILToRocc.scala 37:25]
        bitsBuffer_4 <= io_in_bits; // @[AXILToRocc.scala 37:25]
      end
    end
  end
endmodule
module RoccToAXIL(
  input         clock,
  input         reset,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits,
  output        io_rocc_ready,
  input         io_rocc_valid,
  input  [4:0]  io_rocc_bits_rd,
  input  [63:0] io_rocc_bits_data
);
  reg [63:0] buffer; // @[RoccToAXIL.scala 27:19]
  reg [4:0] rd; // @[RoccToAXIL.scala 29:15]
  wire [95:0] wholePayload = {27'h0,rd,buffer[31:0],buffer[63:32]}; // @[Cat.scala 33:92]
  wire [31:0] beats_0 = wholePayload[31:0]; // @[RoccToAXIL.scala 32:17]
  wire [31:0] beats_1 = wholePayload[63:32]; // @[RoccToAXIL.scala 32:17]
  wire [31:0] beats_2 = wholePayload[95:64]; // @[RoccToAXIL.scala 32:17]
  reg [1:0] beatCounter; // @[RoccToAXIL.scala 34:24]
  reg  state; // @[RoccToAXIL.scala 37:22]
  wire  _io_rocc_ready_T = ~state; // @[RoccToAXIL.scala 40:27]
  wire  _T_1 = io_rocc_ready & io_rocc_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_2 = _T_1 | state; // @[RoccToAXIL.scala 43:26 46:15 37:22]
  wire [31:0] _GEN_5 = 2'h1 == beatCounter ? beats_1 : beats_0; // @[RoccToAXIL.scala 52:{19,19}]
  wire  _T_3 = io_out_ready & io_out_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_7 = beatCounter == 2'h2 ? 1'h0 : state; // @[RoccToAXIL.scala 54:46 55:17 37:22]
  wire [1:0] _beatCounter_T_1 = beatCounter + 2'h1; // @[RoccToAXIL.scala 57:36]
  assign io_out_valid = _io_rocc_ready_T ? 1'h0 : state; // @[RoccToAXIL.scala 38:16 41:17]
  assign io_out_bits = 2'h2 == beatCounter ? beats_2 : _GEN_5; // @[RoccToAXIL.scala 52:{19,19}]
  assign io_rocc_ready = ~state; // @[RoccToAXIL.scala 40:27]
  always @(posedge clock) begin
    if (_io_rocc_ready_T) begin // @[RoccToAXIL.scala 41:17]
      if (_T_1) begin // @[RoccToAXIL.scala 43:26]
        buffer <= io_rocc_bits_data; // @[RoccToAXIL.scala 44:16]
      end
    end
    if (_io_rocc_ready_T) begin // @[RoccToAXIL.scala 41:17]
      if (_T_1) begin // @[RoccToAXIL.scala 43:26]
        rd <= io_rocc_bits_rd; // @[RoccToAXIL.scala 45:12]
      end
    end
    if (_io_rocc_ready_T) begin // @[RoccToAXIL.scala 41:17]
      if (_T_1) begin // @[RoccToAXIL.scala 43:26]
        beatCounter <= 2'h0; // @[RoccToAXIL.scala 47:21]
      end
    end else if (state) begin // @[RoccToAXIL.scala 41:17]
      if (_T_3) begin // @[RoccToAXIL.scala 53:25]
        beatCounter <= _beatCounter_T_1; // @[RoccToAXIL.scala 57:21]
      end
    end
    if (reset) begin // @[RoccToAXIL.scala 37:22]
      state <= 1'h0; // @[RoccToAXIL.scala 37:22]
    end else if (_io_rocc_ready_T) begin // @[RoccToAXIL.scala 41:17]
      state <= _GEN_2;
    end else if (state) begin // @[RoccToAXIL.scala 41:17]
      if (_T_3) begin // @[RoccToAXIL.scala 53:25]
        state <= _GEN_7;
      end
    end
  end
endmodule
module AXILHub(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [15:0] auto_in_aw_bits_id,
  input  [15:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [1:0]  auto_in_aw_bits_burst,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [15:0] auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [15:0] auto_in_ar_bits_id,
  input  [15:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [1:0]  auto_in_ar_bits_burst,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [15:0] auto_in_r_bits_id,
  output [31:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         io_rocc_in_ready,
  output        io_rocc_in_valid,
  output [6:0]  io_rocc_in_bits_inst_funct,
  output [4:0]  io_rocc_in_bits_inst_rs2,
  output [4:0]  io_rocc_in_bits_inst_rs1,
  output [6:0]  io_rocc_in_bits_inst_opcode,
  output [63:0] io_rocc_in_bits_rs1,
  output [63:0] io_rocc_in_bits_rs2,
  output        io_rocc_out_ready,
  input         io_rocc_out_valid,
  input  [4:0]  io_rocc_out_bits_rd,
  input  [63:0] io_rocc_out_bits_data
);
  wire  axil_widget_clock; // @[AXILHub.scala 13:31]
  wire  axil_widget_reset; // @[AXILHub.scala 13:31]
  wire  axil_widget_auto_in_aw_ready; // @[AXILHub.scala 13:31]
  wire  axil_widget_auto_in_aw_valid; // @[AXILHub.scala 13:31]
  wire [15:0] axil_widget_auto_in_aw_bits_id; // @[AXILHub.scala 13:31]
  wire [15:0] axil_widget_auto_in_aw_bits_addr; // @[AXILHub.scala 13:31]
  wire [7:0] axil_widget_auto_in_aw_bits_len; // @[AXILHub.scala 13:31]
  wire [2:0] axil_widget_auto_in_aw_bits_size; // @[AXILHub.scala 13:31]
  wire [1:0] axil_widget_auto_in_aw_bits_burst; // @[AXILHub.scala 13:31]
  wire  axil_widget_auto_in_w_ready; // @[AXILHub.scala 13:31]
  wire  axil_widget_auto_in_w_valid; // @[AXILHub.scala 13:31]
  wire [31:0] axil_widget_auto_in_w_bits_data; // @[AXILHub.scala 13:31]
  wire  axil_widget_auto_in_w_bits_last; // @[AXILHub.scala 13:31]
  wire  axil_widget_auto_in_b_ready; // @[AXILHub.scala 13:31]
  wire  axil_widget_auto_in_b_valid; // @[AXILHub.scala 13:31]
  wire [15:0] axil_widget_auto_in_b_bits_id; // @[AXILHub.scala 13:31]
  wire [1:0] axil_widget_auto_in_b_bits_resp; // @[AXILHub.scala 13:31]
  wire  axil_widget_auto_in_ar_ready; // @[AXILHub.scala 13:31]
  wire  axil_widget_auto_in_ar_valid; // @[AXILHub.scala 13:31]
  wire [15:0] axil_widget_auto_in_ar_bits_id; // @[AXILHub.scala 13:31]
  wire [15:0] axil_widget_auto_in_ar_bits_addr; // @[AXILHub.scala 13:31]
  wire [7:0] axil_widget_auto_in_ar_bits_len; // @[AXILHub.scala 13:31]
  wire [2:0] axil_widget_auto_in_ar_bits_size; // @[AXILHub.scala 13:31]
  wire [1:0] axil_widget_auto_in_ar_bits_burst; // @[AXILHub.scala 13:31]
  wire  axil_widget_auto_in_r_ready; // @[AXILHub.scala 13:31]
  wire  axil_widget_auto_in_r_valid; // @[AXILHub.scala 13:31]
  wire [15:0] axil_widget_auto_in_r_bits_id; // @[AXILHub.scala 13:31]
  wire [31:0] axil_widget_auto_in_r_bits_data; // @[AXILHub.scala 13:31]
  wire [1:0] axil_widget_auto_in_r_bits_resp; // @[AXILHub.scala 13:31]
  wire  axil_widget_auto_in_r_bits_last; // @[AXILHub.scala 13:31]
  wire  axil_widget_io_cmds_ready; // @[AXILHub.scala 13:31]
  wire  axil_widget_io_cmds_valid; // @[AXILHub.scala 13:31]
  wire [31:0] axil_widget_io_cmds_bits; // @[AXILHub.scala 13:31]
  wire  axil_widget_io_resp_ready; // @[AXILHub.scala 13:31]
  wire  axil_widget_io_resp_valid; // @[AXILHub.scala 13:31]
  wire [31:0] axil_widget_io_resp_bits; // @[AXILHub.scala 13:31]
  wire  axil_to_rocc_clock; // @[AXILHub.scala 29:28]
  wire  axil_to_rocc_reset; // @[AXILHub.scala 29:28]
  wire  axil_to_rocc_io_in_ready; // @[AXILHub.scala 29:28]
  wire  axil_to_rocc_io_in_valid; // @[AXILHub.scala 29:28]
  wire [31:0] axil_to_rocc_io_in_bits; // @[AXILHub.scala 29:28]
  wire  axil_to_rocc_io_rocc_ready; // @[AXILHub.scala 29:28]
  wire  axil_to_rocc_io_rocc_valid; // @[AXILHub.scala 29:28]
  wire [6:0] axil_to_rocc_io_rocc_bits_inst_funct; // @[AXILHub.scala 29:28]
  wire [4:0] axil_to_rocc_io_rocc_bits_inst_rs2; // @[AXILHub.scala 29:28]
  wire [4:0] axil_to_rocc_io_rocc_bits_inst_rs1; // @[AXILHub.scala 29:28]
  wire [6:0] axil_to_rocc_io_rocc_bits_inst_opcode; // @[AXILHub.scala 29:28]
  wire [63:0] axil_to_rocc_io_rocc_bits_rs1; // @[AXILHub.scala 29:28]
  wire [63:0] axil_to_rocc_io_rocc_bits_rs2; // @[AXILHub.scala 29:28]
  wire  rocc_to_axil_clock; // @[AXILHub.scala 30:28]
  wire  rocc_to_axil_reset; // @[AXILHub.scala 30:28]
  wire  rocc_to_axil_io_out_ready; // @[AXILHub.scala 30:28]
  wire  rocc_to_axil_io_out_valid; // @[AXILHub.scala 30:28]
  wire [31:0] rocc_to_axil_io_out_bits; // @[AXILHub.scala 30:28]
  wire  rocc_to_axil_io_rocc_ready; // @[AXILHub.scala 30:28]
  wire  rocc_to_axil_io_rocc_valid; // @[AXILHub.scala 30:28]
  wire [4:0] rocc_to_axil_io_rocc_bits_rd; // @[AXILHub.scala 30:28]
  wire [63:0] rocc_to_axil_io_rocc_bits_data; // @[AXILHub.scala 30:28]
  AXILWidget axil_widget ( // @[AXILHub.scala 13:31]
    .clock(axil_widget_clock),
    .reset(axil_widget_reset),
    .auto_in_aw_ready(axil_widget_auto_in_aw_ready),
    .auto_in_aw_valid(axil_widget_auto_in_aw_valid),
    .auto_in_aw_bits_id(axil_widget_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axil_widget_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axil_widget_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axil_widget_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axil_widget_auto_in_aw_bits_burst),
    .auto_in_w_ready(axil_widget_auto_in_w_ready),
    .auto_in_w_valid(axil_widget_auto_in_w_valid),
    .auto_in_w_bits_data(axil_widget_auto_in_w_bits_data),
    .auto_in_w_bits_last(axil_widget_auto_in_w_bits_last),
    .auto_in_b_ready(axil_widget_auto_in_b_ready),
    .auto_in_b_valid(axil_widget_auto_in_b_valid),
    .auto_in_b_bits_id(axil_widget_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axil_widget_auto_in_b_bits_resp),
    .auto_in_ar_ready(axil_widget_auto_in_ar_ready),
    .auto_in_ar_valid(axil_widget_auto_in_ar_valid),
    .auto_in_ar_bits_id(axil_widget_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axil_widget_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axil_widget_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axil_widget_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axil_widget_auto_in_ar_bits_burst),
    .auto_in_r_ready(axil_widget_auto_in_r_ready),
    .auto_in_r_valid(axil_widget_auto_in_r_valid),
    .auto_in_r_bits_id(axil_widget_auto_in_r_bits_id),
    .auto_in_r_bits_data(axil_widget_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axil_widget_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axil_widget_auto_in_r_bits_last),
    .io_cmds_ready(axil_widget_io_cmds_ready),
    .io_cmds_valid(axil_widget_io_cmds_valid),
    .io_cmds_bits(axil_widget_io_cmds_bits),
    .io_resp_ready(axil_widget_io_resp_ready),
    .io_resp_valid(axil_widget_io_resp_valid),
    .io_resp_bits(axil_widget_io_resp_bits)
  );
  AXILToRocc axil_to_rocc ( // @[AXILHub.scala 29:28]
    .clock(axil_to_rocc_clock),
    .reset(axil_to_rocc_reset),
    .io_in_ready(axil_to_rocc_io_in_ready),
    .io_in_valid(axil_to_rocc_io_in_valid),
    .io_in_bits(axil_to_rocc_io_in_bits),
    .io_rocc_ready(axil_to_rocc_io_rocc_ready),
    .io_rocc_valid(axil_to_rocc_io_rocc_valid),
    .io_rocc_bits_inst_funct(axil_to_rocc_io_rocc_bits_inst_funct),
    .io_rocc_bits_inst_rs2(axil_to_rocc_io_rocc_bits_inst_rs2),
    .io_rocc_bits_inst_rs1(axil_to_rocc_io_rocc_bits_inst_rs1),
    .io_rocc_bits_inst_opcode(axil_to_rocc_io_rocc_bits_inst_opcode),
    .io_rocc_bits_rs1(axil_to_rocc_io_rocc_bits_rs1),
    .io_rocc_bits_rs2(axil_to_rocc_io_rocc_bits_rs2)
  );
  RoccToAXIL rocc_to_axil ( // @[AXILHub.scala 30:28]
    .clock(rocc_to_axil_clock),
    .reset(rocc_to_axil_reset),
    .io_out_ready(rocc_to_axil_io_out_ready),
    .io_out_valid(rocc_to_axil_io_out_valid),
    .io_out_bits(rocc_to_axil_io_out_bits),
    .io_rocc_ready(rocc_to_axil_io_rocc_ready),
    .io_rocc_valid(rocc_to_axil_io_rocc_valid),
    .io_rocc_bits_rd(rocc_to_axil_io_rocc_bits_rd),
    .io_rocc_bits_data(rocc_to_axil_io_rocc_bits_data)
  );
  assign auto_in_aw_ready = axil_widget_auto_in_aw_ready; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign auto_in_w_ready = axil_widget_auto_in_w_ready; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign auto_in_b_valid = axil_widget_auto_in_b_valid; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign auto_in_b_bits_id = axil_widget_auto_in_b_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign auto_in_b_bits_resp = axil_widget_auto_in_b_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign auto_in_ar_ready = axil_widget_auto_in_ar_ready; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign auto_in_r_valid = axil_widget_auto_in_r_valid; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign auto_in_r_bits_id = axil_widget_auto_in_r_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign auto_in_r_bits_data = axil_widget_auto_in_r_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign auto_in_r_bits_resp = axil_widget_auto_in_r_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign auto_in_r_bits_last = axil_widget_auto_in_r_bits_last; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign io_rocc_in_valid = axil_to_rocc_io_rocc_valid; // @[AXILHub.scala 35:14]
  assign io_rocc_in_bits_inst_funct = axil_to_rocc_io_rocc_bits_inst_funct; // @[AXILHub.scala 35:14]
  assign io_rocc_in_bits_inst_rs2 = axil_to_rocc_io_rocc_bits_inst_rs2; // @[AXILHub.scala 35:14]
  assign io_rocc_in_bits_inst_rs1 = axil_to_rocc_io_rocc_bits_inst_rs1; // @[AXILHub.scala 35:14]
  assign io_rocc_in_bits_inst_opcode = axil_to_rocc_io_rocc_bits_inst_opcode; // @[AXILHub.scala 35:14]
  assign io_rocc_in_bits_rs1 = axil_to_rocc_io_rocc_bits_rs1; // @[AXILHub.scala 35:14]
  assign io_rocc_in_bits_rs2 = axil_to_rocc_io_rocc_bits_rs2; // @[AXILHub.scala 35:14]
  assign io_rocc_out_ready = rocc_to_axil_io_rocc_ready; // @[AXILHub.scala 33:24]
  assign axil_widget_clock = clock;
  assign axil_widget_reset = reset;
  assign axil_widget_auto_in_aw_valid = auto_in_aw_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axil_widget_auto_in_aw_bits_id = auto_in_aw_bits_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axil_widget_auto_in_aw_bits_addr = auto_in_aw_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axil_widget_auto_in_aw_bits_len = auto_in_aw_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axil_widget_auto_in_aw_bits_size = auto_in_aw_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axil_widget_auto_in_aw_bits_burst = auto_in_aw_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axil_widget_auto_in_w_valid = auto_in_w_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axil_widget_auto_in_w_bits_data = auto_in_w_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axil_widget_auto_in_w_bits_last = auto_in_w_bits_last; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axil_widget_auto_in_b_ready = auto_in_b_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axil_widget_auto_in_ar_valid = auto_in_ar_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axil_widget_auto_in_ar_bits_id = auto_in_ar_bits_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axil_widget_auto_in_ar_bits_addr = auto_in_ar_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axil_widget_auto_in_ar_bits_len = auto_in_ar_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axil_widget_auto_in_ar_bits_size = auto_in_ar_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axil_widget_auto_in_ar_bits_burst = auto_in_ar_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axil_widget_auto_in_r_ready = auto_in_r_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign axil_widget_io_cmds_ready = axil_to_rocc_io_in_ready; // @[AXILHub.scala 34:22]
  assign axil_widget_io_resp_valid = rocc_to_axil_io_out_valid; // @[AXILHub.scala 32:23]
  assign axil_widget_io_resp_bits = rocc_to_axil_io_out_bits; // @[AXILHub.scala 32:23]
  assign axil_to_rocc_clock = clock;
  assign axil_to_rocc_reset = reset;
  assign axil_to_rocc_io_in_valid = axil_widget_io_cmds_valid; // @[AXILHub.scala 34:22]
  assign axil_to_rocc_io_in_bits = axil_widget_io_cmds_bits; // @[AXILHub.scala 34:22]
  assign axil_to_rocc_io_rocc_ready = io_rocc_in_ready; // @[AXILHub.scala 35:14]
  assign rocc_to_axil_clock = clock;
  assign rocc_to_axil_reset = reset;
  assign rocc_to_axil_io_out_ready = axil_widget_io_resp_ready; // @[AXILHub.scala 32:23]
  assign rocc_to_axil_io_rocc_valid = io_rocc_out_valid; // @[AXILHub.scala 33:24]
  assign rocc_to_axil_io_rocc_bits_rd = io_rocc_out_bits_rd; // @[AXILHub.scala 33:24]
  assign rocc_to_axil_io_rocc_bits_data = io_rocc_out_bits_data; // @[AXILHub.scala 33:24]
endmodule
module Queue_182(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [15:0] io_enq_bits_id,
  input  [15:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_len,
  input  [2:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_burst,
  input         io_deq_ready,
  output        io_deq_valid,
  output [15:0] io_deq_bits_id,
  output [15:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_len,
  output [2:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_burst
);
  reg [15:0] ram_id [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [15:0] ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [15:0] ram_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [15:0] ram_addr [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_addr_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_addr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [15:0] ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [15:0] ram_addr_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_addr_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_addr_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_addr_MPORT_en; // @[Decoupled.scala 273:95]
  reg [7:0] ram_len [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_len_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_len_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [7:0] ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [7:0] ram_len_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_len_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_len_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_len_MPORT_en; // @[Decoupled.scala 273:95]
  reg [2:0] ram_size [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [2:0] ram_size_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_burst [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_burst_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_burst_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_burst_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_burst_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_burst_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_burst_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = enq_ptr_value;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_addr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_addr_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = enq_ptr_value;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_len_io_deq_bits_MPORT_en = 1'h1;
  assign ram_len_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_len_io_deq_bits_MPORT_data = ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_len_MPORT_data = io_enq_bits_len;
  assign ram_len_MPORT_addr = enq_ptr_value;
  assign ram_len_MPORT_mask = 1'h1;
  assign ram_len_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = enq_ptr_value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_burst_io_deq_bits_MPORT_en = 1'h1;
  assign ram_burst_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_burst_io_deq_bits_MPORT_data = ram_burst[ram_burst_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_burst_MPORT_data = io_enq_bits_burst;
  assign ram_burst_MPORT_addr = enq_ptr_value;
  assign ram_burst_MPORT_mask = 1'h1;
  assign ram_burst_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_id = ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_addr = ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_len = ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_burst = ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_len_MPORT_en & ram_len_MPORT_mask) begin
      ram_len[ram_len_MPORT_addr] <= ram_len_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_burst_MPORT_en & ram_burst_MPORT_mask) begin
      ram_burst[ram_burst_MPORT_addr] <= ram_burst_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
endmodule
module Queue_183(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] ram_data [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [31:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [31:0] ram_data_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_last [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_last_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_last_io_deq_bits_MPORT_data = ram_last[ram_last_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_last_MPORT_data = io_enq_bits_last;
  assign ram_last_MPORT_addr = enq_ptr_value;
  assign ram_last_MPORT_mask = 1'h1;
  assign ram_last_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_last = ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_last_MPORT_en & ram_last_MPORT_mask) begin
      ram_last[ram_last_MPORT_addr] <= ram_last_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
endmodule
module Queue_184(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [15:0] io_enq_bits_id,
  input  [1:0]  io_enq_bits_resp,
  input         io_deq_ready,
  output        io_deq_valid,
  output [15:0] io_deq_bits_id,
  output [1:0]  io_deq_bits_resp
);
  reg [15:0] ram_id [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [15:0] ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [15:0] ram_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_resp [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_resp_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_resp_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_resp_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = enq_ptr_value;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_resp_io_deq_bits_MPORT_en = 1'h1;
  assign ram_resp_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_resp_io_deq_bits_MPORT_data = ram_resp[ram_resp_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_resp_MPORT_data = io_enq_bits_resp;
  assign ram_resp_MPORT_addr = enq_ptr_value;
  assign ram_resp_MPORT_mask = 1'h1;
  assign ram_resp_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_id = ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_resp = ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_resp_MPORT_en & ram_resp_MPORT_mask) begin
      ram_resp[ram_resp_MPORT_addr] <= ram_resp_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
endmodule
module Queue_186(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [15:0] io_enq_bits_id,
  input  [31:0] io_enq_bits_data,
  input  [1:0]  io_enq_bits_resp,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [15:0] io_deq_bits_id,
  output [31:0] io_deq_bits_data,
  output [1:0]  io_deq_bits_resp,
  output        io_deq_bits_last
);
  reg [15:0] ram_id [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [15:0] ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [15:0] ram_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [31:0] ram_data [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [31:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [31:0] ram_data_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_resp [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_resp_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_resp_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_resp_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_resp_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_last [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_last_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = enq_ptr_value;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_resp_io_deq_bits_MPORT_en = 1'h1;
  assign ram_resp_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_resp_io_deq_bits_MPORT_data = ram_resp[ram_resp_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_resp_MPORT_data = io_enq_bits_resp;
  assign ram_resp_MPORT_addr = enq_ptr_value;
  assign ram_resp_MPORT_mask = 1'h1;
  assign ram_resp_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_last_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_last_io_deq_bits_MPORT_data = ram_last[ram_last_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_last_MPORT_data = io_enq_bits_last;
  assign ram_last_MPORT_addr = enq_ptr_value;
  assign ram_last_MPORT_mask = 1'h1;
  assign ram_last_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_id = ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_resp = ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_last = ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_resp_MPORT_en & ram_resp_MPORT_mask) begin
      ram_resp[ram_resp_MPORT_addr] <= ram_resp_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_last_MPORT_en & ram_last_MPORT_mask) begin
      ram_last[ram_last_MPORT_addr] <= ram_last_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
endmodule
module AXI4Buffer_6(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [15:0] auto_in_aw_bits_id,
  input  [15:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [1:0]  auto_in_aw_bits_burst,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [15:0] auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [15:0] auto_in_ar_bits_id,
  input  [15:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [1:0]  auto_in_ar_bits_burst,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [15:0] auto_in_r_bits_id,
  output [31:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output [15:0] auto_out_aw_bits_id,
  output [15:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  output [1:0]  auto_out_aw_bits_burst,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [31:0] auto_out_w_bits_data,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [15:0] auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output [15:0] auto_out_ar_bits_id,
  output [15:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output [1:0]  auto_out_ar_bits_burst,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [15:0] auto_out_r_bits_id,
  input  [31:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input         auto_out_r_bits_last
);
  wire  x1_aw_deq_clock; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_reset; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [15:0] x1_aw_deq_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire [15:0] x1_aw_deq_io_enq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] x1_aw_deq_io_enq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] x1_aw_deq_io_enq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] x1_aw_deq_io_enq_bits_burst; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  x1_aw_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [15:0] x1_aw_deq_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [15:0] x1_aw_deq_io_deq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] x1_aw_deq_io_deq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] x1_aw_deq_io_deq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] x1_aw_deq_io_deq_bits_burst; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_clock; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_reset; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [31:0] x1_w_deq_io_enq_bits_data; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_enq_bits_last; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [31:0] x1_w_deq_io_deq_bits_data; // @[Decoupled.scala 375:21]
  wire  x1_w_deq_io_deq_bits_last; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_clock; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_reset; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [15:0] bundleIn_0_b_deq_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire [1:0] bundleIn_0_b_deq_io_enq_bits_resp; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_b_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [15:0] bundleIn_0_b_deq_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [1:0] bundleIn_0_b_deq_io_deq_bits_resp; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_clock; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_reset; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [15:0] x1_ar_deq_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire [15:0] x1_ar_deq_io_enq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] x1_ar_deq_io_enq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] x1_ar_deq_io_enq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] x1_ar_deq_io_enq_bits_burst; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  x1_ar_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [15:0] x1_ar_deq_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [15:0] x1_ar_deq_io_deq_bits_addr; // @[Decoupled.scala 375:21]
  wire [7:0] x1_ar_deq_io_deq_bits_len; // @[Decoupled.scala 375:21]
  wire [2:0] x1_ar_deq_io_deq_bits_size; // @[Decoupled.scala 375:21]
  wire [1:0] x1_ar_deq_io_deq_bits_burst; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_clock; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_reset; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_enq_valid; // @[Decoupled.scala 375:21]
  wire [15:0] bundleIn_0_r_deq_io_enq_bits_id; // @[Decoupled.scala 375:21]
  wire [31:0] bundleIn_0_r_deq_io_enq_bits_data; // @[Decoupled.scala 375:21]
  wire [1:0] bundleIn_0_r_deq_io_enq_bits_resp; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_enq_bits_last; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_deq_valid; // @[Decoupled.scala 375:21]
  wire [15:0] bundleIn_0_r_deq_io_deq_bits_id; // @[Decoupled.scala 375:21]
  wire [31:0] bundleIn_0_r_deq_io_deq_bits_data; // @[Decoupled.scala 375:21]
  wire [1:0] bundleIn_0_r_deq_io_deq_bits_resp; // @[Decoupled.scala 375:21]
  wire  bundleIn_0_r_deq_io_deq_bits_last; // @[Decoupled.scala 375:21]
  Queue_182 x1_aw_deq ( // @[Decoupled.scala 375:21]
    .clock(x1_aw_deq_clock),
    .reset(x1_aw_deq_reset),
    .io_enq_ready(x1_aw_deq_io_enq_ready),
    .io_enq_valid(x1_aw_deq_io_enq_valid),
    .io_enq_bits_id(x1_aw_deq_io_enq_bits_id),
    .io_enq_bits_addr(x1_aw_deq_io_enq_bits_addr),
    .io_enq_bits_len(x1_aw_deq_io_enq_bits_len),
    .io_enq_bits_size(x1_aw_deq_io_enq_bits_size),
    .io_enq_bits_burst(x1_aw_deq_io_enq_bits_burst),
    .io_deq_ready(x1_aw_deq_io_deq_ready),
    .io_deq_valid(x1_aw_deq_io_deq_valid),
    .io_deq_bits_id(x1_aw_deq_io_deq_bits_id),
    .io_deq_bits_addr(x1_aw_deq_io_deq_bits_addr),
    .io_deq_bits_len(x1_aw_deq_io_deq_bits_len),
    .io_deq_bits_size(x1_aw_deq_io_deq_bits_size),
    .io_deq_bits_burst(x1_aw_deq_io_deq_bits_burst)
  );
  Queue_183 x1_w_deq ( // @[Decoupled.scala 375:21]
    .clock(x1_w_deq_clock),
    .reset(x1_w_deq_reset),
    .io_enq_ready(x1_w_deq_io_enq_ready),
    .io_enq_valid(x1_w_deq_io_enq_valid),
    .io_enq_bits_data(x1_w_deq_io_enq_bits_data),
    .io_enq_bits_last(x1_w_deq_io_enq_bits_last),
    .io_deq_ready(x1_w_deq_io_deq_ready),
    .io_deq_valid(x1_w_deq_io_deq_valid),
    .io_deq_bits_data(x1_w_deq_io_deq_bits_data),
    .io_deq_bits_last(x1_w_deq_io_deq_bits_last)
  );
  Queue_184 bundleIn_0_b_deq ( // @[Decoupled.scala 375:21]
    .clock(bundleIn_0_b_deq_clock),
    .reset(bundleIn_0_b_deq_reset),
    .io_enq_ready(bundleIn_0_b_deq_io_enq_ready),
    .io_enq_valid(bundleIn_0_b_deq_io_enq_valid),
    .io_enq_bits_id(bundleIn_0_b_deq_io_enq_bits_id),
    .io_enq_bits_resp(bundleIn_0_b_deq_io_enq_bits_resp),
    .io_deq_ready(bundleIn_0_b_deq_io_deq_ready),
    .io_deq_valid(bundleIn_0_b_deq_io_deq_valid),
    .io_deq_bits_id(bundleIn_0_b_deq_io_deq_bits_id),
    .io_deq_bits_resp(bundleIn_0_b_deq_io_deq_bits_resp)
  );
  Queue_182 x1_ar_deq ( // @[Decoupled.scala 375:21]
    .clock(x1_ar_deq_clock),
    .reset(x1_ar_deq_reset),
    .io_enq_ready(x1_ar_deq_io_enq_ready),
    .io_enq_valid(x1_ar_deq_io_enq_valid),
    .io_enq_bits_id(x1_ar_deq_io_enq_bits_id),
    .io_enq_bits_addr(x1_ar_deq_io_enq_bits_addr),
    .io_enq_bits_len(x1_ar_deq_io_enq_bits_len),
    .io_enq_bits_size(x1_ar_deq_io_enq_bits_size),
    .io_enq_bits_burst(x1_ar_deq_io_enq_bits_burst),
    .io_deq_ready(x1_ar_deq_io_deq_ready),
    .io_deq_valid(x1_ar_deq_io_deq_valid),
    .io_deq_bits_id(x1_ar_deq_io_deq_bits_id),
    .io_deq_bits_addr(x1_ar_deq_io_deq_bits_addr),
    .io_deq_bits_len(x1_ar_deq_io_deq_bits_len),
    .io_deq_bits_size(x1_ar_deq_io_deq_bits_size),
    .io_deq_bits_burst(x1_ar_deq_io_deq_bits_burst)
  );
  Queue_186 bundleIn_0_r_deq ( // @[Decoupled.scala 375:21]
    .clock(bundleIn_0_r_deq_clock),
    .reset(bundleIn_0_r_deq_reset),
    .io_enq_ready(bundleIn_0_r_deq_io_enq_ready),
    .io_enq_valid(bundleIn_0_r_deq_io_enq_valid),
    .io_enq_bits_id(bundleIn_0_r_deq_io_enq_bits_id),
    .io_enq_bits_data(bundleIn_0_r_deq_io_enq_bits_data),
    .io_enq_bits_resp(bundleIn_0_r_deq_io_enq_bits_resp),
    .io_enq_bits_last(bundleIn_0_r_deq_io_enq_bits_last),
    .io_deq_ready(bundleIn_0_r_deq_io_deq_ready),
    .io_deq_valid(bundleIn_0_r_deq_io_deq_valid),
    .io_deq_bits_id(bundleIn_0_r_deq_io_deq_bits_id),
    .io_deq_bits_data(bundleIn_0_r_deq_io_deq_bits_data),
    .io_deq_bits_resp(bundleIn_0_r_deq_io_deq_bits_resp),
    .io_deq_bits_last(bundleIn_0_r_deq_io_deq_bits_last)
  );
  assign auto_in_aw_ready = x1_aw_deq_io_enq_ready; // @[Nodes.scala 1215:84 Decoupled.scala 379:17]
  assign auto_in_w_ready = x1_w_deq_io_enq_ready; // @[Nodes.scala 1215:84 Decoupled.scala 379:17]
  assign auto_in_b_valid = bundleIn_0_b_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_in_b_bits_id = bundleIn_0_b_deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_b_bits_resp = bundleIn_0_b_deq_io_deq_bits_resp; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_ar_ready = x1_ar_deq_io_enq_ready; // @[Nodes.scala 1215:84 Decoupled.scala 379:17]
  assign auto_in_r_valid = bundleIn_0_r_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_in_r_bits_id = bundleIn_0_r_deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_r_bits_data = bundleIn_0_r_deq_io_deq_bits_data; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_r_bits_resp = bundleIn_0_r_deq_io_deq_bits_resp; // @[Decoupled.scala 414:19 415:14]
  assign auto_in_r_bits_last = bundleIn_0_r_deq_io_deq_bits_last; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_valid = x1_aw_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_out_aw_bits_id = x1_aw_deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_addr = x1_aw_deq_io_deq_bits_addr; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_len = x1_aw_deq_io_deq_bits_len; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_size = x1_aw_deq_io_deq_bits_size; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_aw_bits_burst = x1_aw_deq_io_deq_bits_burst; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_w_valid = x1_w_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_out_w_bits_data = x1_w_deq_io_deq_bits_data; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_w_bits_last = x1_w_deq_io_deq_bits_last; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_b_ready = bundleIn_0_b_deq_io_enq_ready; // @[Nodes.scala 1212:84 Decoupled.scala 379:17]
  assign auto_out_ar_valid = x1_ar_deq_io_deq_valid; // @[Decoupled.scala 414:19 416:15]
  assign auto_out_ar_bits_id = x1_ar_deq_io_deq_bits_id; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_addr = x1_ar_deq_io_deq_bits_addr; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_len = x1_ar_deq_io_deq_bits_len; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_size = x1_ar_deq_io_deq_bits_size; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_ar_bits_burst = x1_ar_deq_io_deq_bits_burst; // @[Decoupled.scala 414:19 415:14]
  assign auto_out_r_ready = bundleIn_0_r_deq_io_enq_ready; // @[Nodes.scala 1212:84 Decoupled.scala 379:17]
  assign x1_aw_deq_clock = clock;
  assign x1_aw_deq_reset = reset;
  assign x1_aw_deq_io_enq_valid = auto_in_aw_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_id = auto_in_aw_bits_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_addr = auto_in_aw_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_len = auto_in_aw_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_size = auto_in_aw_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_enq_bits_burst = auto_in_aw_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_aw_deq_io_deq_ready = auto_out_aw_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign x1_w_deq_clock = clock;
  assign x1_w_deq_reset = reset;
  assign x1_w_deq_io_enq_valid = auto_in_w_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_w_deq_io_enq_bits_data = auto_in_w_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_w_deq_io_enq_bits_last = auto_in_w_bits_last; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_w_deq_io_deq_ready = auto_out_w_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_b_deq_clock = clock;
  assign bundleIn_0_b_deq_reset = reset;
  assign bundleIn_0_b_deq_io_enq_valid = auto_out_b_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_b_deq_io_enq_bits_id = auto_out_b_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_b_deq_io_enq_bits_resp = auto_out_b_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_b_deq_io_deq_ready = auto_in_b_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_clock = clock;
  assign x1_ar_deq_reset = reset;
  assign x1_ar_deq_io_enq_valid = auto_in_ar_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_id = auto_in_ar_bits_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_addr = auto_in_ar_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_len = auto_in_ar_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_size = auto_in_ar_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_enq_bits_burst = auto_in_ar_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign x1_ar_deq_io_deq_ready = auto_out_ar_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_clock = clock;
  assign bundleIn_0_r_deq_reset = reset;
  assign bundleIn_0_r_deq_io_enq_valid = auto_out_r_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_enq_bits_id = auto_out_r_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_enq_bits_data = auto_out_r_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_enq_bits_resp = auto_out_r_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_enq_bits_last = auto_out_r_bits_last; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign bundleIn_0_r_deq_io_deq_ready = auto_in_r_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
endmodule
module ComposerTop(
  input          clock,
  input          reset,
  input  [15:0]  S00_AXI_awid,
  input  [15:0]  S00_AXI_awaddr,
  input  [7:0]   S00_AXI_awlen,
  input  [2:0]   S00_AXI_awsize,
  input  [1:0]   S00_AXI_awburst,
  input          S00_AXI_awlock,
  input  [3:0]   S00_AXI_awcache,
  input  [2:0]   S00_AXI_awprot,
  input  [3:0]   S00_AXI_awregion,
  input  [3:0]   S00_AXI_awqos,
  input          S00_AXI_awvalid,
  output         S00_AXI_awready,
  input  [31:0]  S00_AXI_wdata,
  input  [3:0]   S00_AXI_wstrb,
  input          S00_AXI_wlast,
  input          S00_AXI_wvalid,
  output         S00_AXI_wready,
  output [15:0]  S00_AXI_bid,
  output [1:0]   S00_AXI_bresp,
  output         S00_AXI_bvalid,
  input          S00_AXI_bready,
  input  [15:0]  S00_AXI_arid,
  input  [15:0]  S00_AXI_araddr,
  input  [7:0]   S00_AXI_arlen,
  input  [2:0]   S00_AXI_arsize,
  input  [1:0]   S00_AXI_arburst,
  input          S00_AXI_arlock,
  input  [3:0]   S00_AXI_arcache,
  input  [2:0]   S00_AXI_arprot,
  input  [3:0]   S00_AXI_arregion,
  input  [3:0]   S00_AXI_arqos,
  input          S00_AXI_arvalid,
  output         S00_AXI_arready,
  output [15:0]  S00_AXI_rid,
  output [31:0]  S00_AXI_rdata,
  output [1:0]   S00_AXI_rresp,
  output         S00_AXI_rlast,
  output         S00_AXI_rvalid,
  input          S00_AXI_rready,
  output [5:0]   M00_AXI_awid,
  output [33:0]  M00_AXI_awaddr,
  output [7:0]   M00_AXI_awlen,
  output [2:0]   M00_AXI_awsize,
  output [1:0]   M00_AXI_awburst,
  output         M00_AXI_awlock,
  output [3:0]   M00_AXI_awcache,
  output [2:0]   M00_AXI_awprot,
  output [3:0]   M00_AXI_awregion,
  output [3:0]   M00_AXI_awqos,
  output         M00_AXI_awvalid,
  input          M00_AXI_awready,
  output [511:0] M00_AXI_wdata,
  output [63:0]  M00_AXI_wstrb,
  output         M00_AXI_wlast,
  output         M00_AXI_wvalid,
  input          M00_AXI_wready,
  input  [5:0]   M00_AXI_bid,
  input  [1:0]   M00_AXI_bresp,
  input          M00_AXI_bvalid,
  output         M00_AXI_bready,
  output [5:0]   M00_AXI_arid,
  output [33:0]  M00_AXI_araddr,
  output [7:0]   M00_AXI_arlen,
  output [2:0]   M00_AXI_arsize,
  output [1:0]   M00_AXI_arburst,
  output         M00_AXI_arlock,
  output [3:0]   M00_AXI_arcache,
  output [2:0]   M00_AXI_arprot,
  output [3:0]   M00_AXI_arregion,
  output [3:0]   M00_AXI_arqos,
  output         M00_AXI_arvalid,
  input          M00_AXI_arready,
  input  [5:0]   M00_AXI_rid,
  input  [511:0] M00_AXI_rdata,
  input  [1:0]   M00_AXI_rresp,
  input          M00_AXI_rlast,
  input          M00_AXI_rvalid,
  output         M00_AXI_rready,
  input  [5:0]   dma_awid,
  input  [33:0]  dma_awaddr,
  input  [7:0]   dma_awlen,
  input  [2:0]   dma_awsize,
  input  [1:0]   dma_awburst,
  input          dma_awlock,
  input  [3:0]   dma_awcache,
  input  [2:0]   dma_awprot,
  input  [3:0]   dma_awregion,
  input  [3:0]   dma_awqos,
  input          dma_awvalid,
  output         dma_awready,
  input  [511:0] dma_wdata,
  input  [63:0]  dma_wstrb,
  input          dma_wlast,
  input          dma_wvalid,
  output         dma_wready,
  output [5:0]   dma_bid,
  output [1:0]   dma_bresp,
  output         dma_bvalid,
  input          dma_bready,
  input  [5:0]   dma_arid,
  input  [33:0]  dma_araddr,
  input  [7:0]   dma_arlen,
  input  [2:0]   dma_arsize,
  input  [1:0]   dma_arburst,
  input          dma_arlock,
  input  [3:0]   dma_arcache,
  input  [2:0]   dma_arprot,
  input  [3:0]   dma_arregion,
  input  [3:0]   dma_arqos,
  input          dma_arvalid,
  output         dma_arready,
  output [5:0]   dma_rid,
  output [511:0] dma_rdata,
  output [1:0]   dma_rresp,
  output         dma_rlast,
  output         dma_rvalid,
  input          dma_rready
);
  wire  acc_clock; // @[ComposerTop.scala 80:23]
  wire  acc_reset; // @[ComposerTop.scala 80:23]
  wire  acc_auto_mem_out_a_ready; // @[ComposerTop.scala 80:23]
  wire  acc_auto_mem_out_a_valid; // @[ComposerTop.scala 80:23]
  wire [2:0] acc_auto_mem_out_a_bits_opcode; // @[ComposerTop.scala 80:23]
  wire [2:0] acc_auto_mem_out_a_bits_size; // @[ComposerTop.scala 80:23]
  wire [6:0] acc_auto_mem_out_a_bits_source; // @[ComposerTop.scala 80:23]
  wire [33:0] acc_auto_mem_out_a_bits_address; // @[ComposerTop.scala 80:23]
  wire [63:0] acc_auto_mem_out_a_bits_mask; // @[ComposerTop.scala 80:23]
  wire [511:0] acc_auto_mem_out_a_bits_data; // @[ComposerTop.scala 80:23]
  wire  acc_auto_mem_out_d_ready; // @[ComposerTop.scala 80:23]
  wire  acc_auto_mem_out_d_valid; // @[ComposerTop.scala 80:23]
  wire [6:0] acc_auto_mem_out_d_bits_source; // @[ComposerTop.scala 80:23]
  wire [511:0] acc_auto_mem_out_d_bits_data; // @[ComposerTop.scala 80:23]
  wire  acc_io_cmd_ready; // @[ComposerTop.scala 80:23]
  wire  acc_io_cmd_valid; // @[ComposerTop.scala 80:23]
  wire [6:0] acc_io_cmd_bits_inst_funct; // @[ComposerTop.scala 80:23]
  wire [4:0] acc_io_cmd_bits_inst_rs2; // @[ComposerTop.scala 80:23]
  wire [4:0] acc_io_cmd_bits_inst_rs1; // @[ComposerTop.scala 80:23]
  wire [6:0] acc_io_cmd_bits_inst_opcode; // @[ComposerTop.scala 80:23]
  wire [63:0] acc_io_cmd_bits_rs1; // @[ComposerTop.scala 80:23]
  wire [63:0] acc_io_cmd_bits_rs2; // @[ComposerTop.scala 80:23]
  wire  acc_io_resp_ready; // @[ComposerTop.scala 80:23]
  wire  acc_io_resp_valid; // @[ComposerTop.scala 80:23]
  wire [4:0] acc_io_resp_bits_rd; // @[ComposerTop.scala 80:23]
  wire [63:0] acc_io_resp_bits_data; // @[ComposerTop.scala 80:23]
  wire  axi4buf_clock; // @[Buffer.scala 63:29]
  wire  axi4buf_reset; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_in_aw_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_in_aw_valid; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_auto_in_aw_bits_id; // @[Buffer.scala 63:29]
  wire [33:0] axi4buf_auto_in_aw_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_auto_in_aw_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_auto_in_aw_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_auto_in_aw_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_in_aw_bits_lock; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_auto_in_aw_bits_cache; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_auto_in_aw_bits_prot; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_auto_in_aw_bits_qos; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_auto_in_aw_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_in_w_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_in_w_valid; // @[Buffer.scala 63:29]
  wire [511:0] axi4buf_auto_in_w_bits_data; // @[Buffer.scala 63:29]
  wire [63:0] axi4buf_auto_in_w_bits_strb; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_in_w_bits_last; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_in_b_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_in_b_valid; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_auto_in_b_bits_id; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_auto_in_b_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_in_ar_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_in_ar_valid; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_auto_in_ar_bits_id; // @[Buffer.scala 63:29]
  wire [33:0] axi4buf_auto_in_ar_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_auto_in_ar_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_auto_in_ar_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_auto_in_ar_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_in_ar_bits_lock; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_auto_in_ar_bits_cache; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_auto_in_ar_bits_prot; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_auto_in_ar_bits_qos; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_auto_in_ar_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_in_r_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_in_r_valid; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_auto_in_r_bits_id; // @[Buffer.scala 63:29]
  wire [511:0] axi4buf_auto_in_r_bits_data; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_auto_in_r_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_in_r_bits_last; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_out_aw_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_out_aw_valid; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_auto_out_aw_bits_id; // @[Buffer.scala 63:29]
  wire [33:0] axi4buf_auto_out_aw_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_auto_out_aw_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_auto_out_aw_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_auto_out_aw_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_out_aw_bits_lock; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_auto_out_aw_bits_cache; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_auto_out_aw_bits_prot; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_auto_out_aw_bits_qos; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_auto_out_aw_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_out_w_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_out_w_valid; // @[Buffer.scala 63:29]
  wire [511:0] axi4buf_auto_out_w_bits_data; // @[Buffer.scala 63:29]
  wire [63:0] axi4buf_auto_out_w_bits_strb; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_out_w_bits_last; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_out_b_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_out_b_valid; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_auto_out_b_bits_id; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_auto_out_b_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_out_ar_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_out_ar_valid; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_auto_out_ar_bits_id; // @[Buffer.scala 63:29]
  wire [33:0] axi4buf_auto_out_ar_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_auto_out_ar_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_auto_out_ar_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_auto_out_ar_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_out_ar_bits_lock; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_auto_out_ar_bits_cache; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_auto_out_ar_bits_prot; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_auto_out_ar_bits_qos; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_auto_out_ar_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_out_r_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_out_r_valid; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_auto_out_r_bits_id; // @[Buffer.scala 63:29]
  wire [511:0] axi4buf_auto_out_r_bits_data; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_auto_out_r_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire  axi4buf_auto_out_r_bits_last; // @[Buffer.scala 63:29]
  wire  axi4buf_1_clock; // @[Buffer.scala 63:29]
  wire  axi4buf_1_reset; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_in_aw_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_in_aw_valid; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_1_auto_in_aw_bits_id; // @[Buffer.scala 63:29]
  wire [33:0] axi4buf_1_auto_in_aw_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_1_auto_in_aw_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_1_auto_in_aw_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_1_auto_in_aw_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_in_aw_bits_lock; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_1_auto_in_aw_bits_cache; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_1_auto_in_aw_bits_prot; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_1_auto_in_aw_bits_qos; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_1_auto_in_aw_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_in_w_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_in_w_valid; // @[Buffer.scala 63:29]
  wire [511:0] axi4buf_1_auto_in_w_bits_data; // @[Buffer.scala 63:29]
  wire [63:0] axi4buf_1_auto_in_w_bits_strb; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_in_w_bits_last; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_in_b_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_in_b_valid; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_1_auto_in_b_bits_id; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_1_auto_in_b_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_in_ar_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_in_ar_valid; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_1_auto_in_ar_bits_id; // @[Buffer.scala 63:29]
  wire [33:0] axi4buf_1_auto_in_ar_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_1_auto_in_ar_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_1_auto_in_ar_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_1_auto_in_ar_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_in_ar_bits_lock; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_1_auto_in_ar_bits_cache; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_1_auto_in_ar_bits_prot; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_1_auto_in_ar_bits_qos; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_1_auto_in_ar_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_in_r_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_in_r_valid; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_1_auto_in_r_bits_id; // @[Buffer.scala 63:29]
  wire [511:0] axi4buf_1_auto_in_r_bits_data; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_1_auto_in_r_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_in_r_bits_last; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_out_aw_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_out_aw_valid; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_1_auto_out_aw_bits_id; // @[Buffer.scala 63:29]
  wire [33:0] axi4buf_1_auto_out_aw_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_1_auto_out_aw_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_1_auto_out_aw_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_1_auto_out_aw_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_out_aw_bits_lock; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_1_auto_out_aw_bits_cache; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_1_auto_out_aw_bits_prot; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_1_auto_out_aw_bits_qos; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_1_auto_out_aw_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_out_w_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_out_w_valid; // @[Buffer.scala 63:29]
  wire [511:0] axi4buf_1_auto_out_w_bits_data; // @[Buffer.scala 63:29]
  wire [63:0] axi4buf_1_auto_out_w_bits_strb; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_out_w_bits_last; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_out_b_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_out_b_valid; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_1_auto_out_b_bits_id; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_1_auto_out_b_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_out_ar_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_out_ar_valid; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_1_auto_out_ar_bits_id; // @[Buffer.scala 63:29]
  wire [33:0] axi4buf_1_auto_out_ar_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_1_auto_out_ar_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_1_auto_out_ar_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_1_auto_out_ar_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_out_ar_bits_lock; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_1_auto_out_ar_bits_cache; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_1_auto_out_ar_bits_prot; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_1_auto_out_ar_bits_qos; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_1_auto_out_ar_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_out_r_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_out_r_valid; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_1_auto_out_r_bits_id; // @[Buffer.scala 63:29]
  wire [511:0] axi4buf_1_auto_out_r_bits_data; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_1_auto_out_r_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire  axi4buf_1_auto_out_r_bits_last; // @[Buffer.scala 63:29]
  wire  tl2axi4_clock; // @[ToAXI4.scala 286:29]
  wire  tl2axi4_reset; // @[ToAXI4.scala 286:29]
  wire  tl2axi4_auto_in_a_ready; // @[ToAXI4.scala 286:29]
  wire  tl2axi4_auto_in_a_valid; // @[ToAXI4.scala 286:29]
  wire [2:0] tl2axi4_auto_in_a_bits_opcode; // @[ToAXI4.scala 286:29]
  wire [2:0] tl2axi4_auto_in_a_bits_size; // @[ToAXI4.scala 286:29]
  wire [6:0] tl2axi4_auto_in_a_bits_source; // @[ToAXI4.scala 286:29]
  wire [33:0] tl2axi4_auto_in_a_bits_address; // @[ToAXI4.scala 286:29]
  wire [63:0] tl2axi4_auto_in_a_bits_mask; // @[ToAXI4.scala 286:29]
  wire [511:0] tl2axi4_auto_in_a_bits_data; // @[ToAXI4.scala 286:29]
  wire  tl2axi4_auto_in_d_ready; // @[ToAXI4.scala 286:29]
  wire  tl2axi4_auto_in_d_valid; // @[ToAXI4.scala 286:29]
  wire [6:0] tl2axi4_auto_in_d_bits_source; // @[ToAXI4.scala 286:29]
  wire [511:0] tl2axi4_auto_in_d_bits_data; // @[ToAXI4.scala 286:29]
  wire  tl2axi4_auto_out_aw_ready; // @[ToAXI4.scala 286:29]
  wire  tl2axi4_auto_out_aw_valid; // @[ToAXI4.scala 286:29]
  wire [6:0] tl2axi4_auto_out_aw_bits_id; // @[ToAXI4.scala 286:29]
  wire [33:0] tl2axi4_auto_out_aw_bits_addr; // @[ToAXI4.scala 286:29]
  wire [7:0] tl2axi4_auto_out_aw_bits_len; // @[ToAXI4.scala 286:29]
  wire [2:0] tl2axi4_auto_out_aw_bits_size; // @[ToAXI4.scala 286:29]
  wire [1:0] tl2axi4_auto_out_aw_bits_burst; // @[ToAXI4.scala 286:29]
  wire  tl2axi4_auto_out_aw_bits_lock; // @[ToAXI4.scala 286:29]
  wire [3:0] tl2axi4_auto_out_aw_bits_cache; // @[ToAXI4.scala 286:29]
  wire [2:0] tl2axi4_auto_out_aw_bits_prot; // @[ToAXI4.scala 286:29]
  wire [3:0] tl2axi4_auto_out_aw_bits_qos; // @[ToAXI4.scala 286:29]
  wire [6:0] tl2axi4_auto_out_aw_bits_echo_tl_state_source; // @[ToAXI4.scala 286:29]
  wire  tl2axi4_auto_out_w_ready; // @[ToAXI4.scala 286:29]
  wire  tl2axi4_auto_out_w_valid; // @[ToAXI4.scala 286:29]
  wire [511:0] tl2axi4_auto_out_w_bits_data; // @[ToAXI4.scala 286:29]
  wire [63:0] tl2axi4_auto_out_w_bits_strb; // @[ToAXI4.scala 286:29]
  wire  tl2axi4_auto_out_w_bits_last; // @[ToAXI4.scala 286:29]
  wire  tl2axi4_auto_out_b_ready; // @[ToAXI4.scala 286:29]
  wire  tl2axi4_auto_out_b_valid; // @[ToAXI4.scala 286:29]
  wire [6:0] tl2axi4_auto_out_b_bits_id; // @[ToAXI4.scala 286:29]
  wire [6:0] tl2axi4_auto_out_b_bits_echo_tl_state_source; // @[ToAXI4.scala 286:29]
  wire  tl2axi4_auto_out_ar_ready; // @[ToAXI4.scala 286:29]
  wire  tl2axi4_auto_out_ar_valid; // @[ToAXI4.scala 286:29]
  wire [6:0] tl2axi4_auto_out_ar_bits_id; // @[ToAXI4.scala 286:29]
  wire [33:0] tl2axi4_auto_out_ar_bits_addr; // @[ToAXI4.scala 286:29]
  wire [7:0] tl2axi4_auto_out_ar_bits_len; // @[ToAXI4.scala 286:29]
  wire [2:0] tl2axi4_auto_out_ar_bits_size; // @[ToAXI4.scala 286:29]
  wire [1:0] tl2axi4_auto_out_ar_bits_burst; // @[ToAXI4.scala 286:29]
  wire  tl2axi4_auto_out_ar_bits_lock; // @[ToAXI4.scala 286:29]
  wire [3:0] tl2axi4_auto_out_ar_bits_cache; // @[ToAXI4.scala 286:29]
  wire [2:0] tl2axi4_auto_out_ar_bits_prot; // @[ToAXI4.scala 286:29]
  wire [3:0] tl2axi4_auto_out_ar_bits_qos; // @[ToAXI4.scala 286:29]
  wire [6:0] tl2axi4_auto_out_ar_bits_echo_tl_state_source; // @[ToAXI4.scala 286:29]
  wire  tl2axi4_auto_out_r_ready; // @[ToAXI4.scala 286:29]
  wire  tl2axi4_auto_out_r_valid; // @[ToAXI4.scala 286:29]
  wire [6:0] tl2axi4_auto_out_r_bits_id; // @[ToAXI4.scala 286:29]
  wire [511:0] tl2axi4_auto_out_r_bits_data; // @[ToAXI4.scala 286:29]
  wire [6:0] tl2axi4_auto_out_r_bits_echo_tl_state_source; // @[ToAXI4.scala 286:29]
  wire  tl2axi4_auto_out_r_bits_last; // @[ToAXI4.scala 286:29]
  wire  axi4xbar_clock; // @[Xbar.scala 231:30]
  wire  axi4xbar_reset; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_1_aw_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_1_aw_valid; // @[Xbar.scala 231:30]
  wire [5:0] axi4xbar_auto_in_1_aw_bits_id; // @[Xbar.scala 231:30]
  wire [33:0] axi4xbar_auto_in_1_aw_bits_addr; // @[Xbar.scala 231:30]
  wire [7:0] axi4xbar_auto_in_1_aw_bits_len; // @[Xbar.scala 231:30]
  wire [2:0] axi4xbar_auto_in_1_aw_bits_size; // @[Xbar.scala 231:30]
  wire [1:0] axi4xbar_auto_in_1_aw_bits_burst; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_1_aw_bits_lock; // @[Xbar.scala 231:30]
  wire [3:0] axi4xbar_auto_in_1_aw_bits_cache; // @[Xbar.scala 231:30]
  wire [2:0] axi4xbar_auto_in_1_aw_bits_prot; // @[Xbar.scala 231:30]
  wire [3:0] axi4xbar_auto_in_1_aw_bits_qos; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_1_w_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_1_w_valid; // @[Xbar.scala 231:30]
  wire [511:0] axi4xbar_auto_in_1_w_bits_data; // @[Xbar.scala 231:30]
  wire [63:0] axi4xbar_auto_in_1_w_bits_strb; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_1_w_bits_last; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_1_b_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_1_b_valid; // @[Xbar.scala 231:30]
  wire [5:0] axi4xbar_auto_in_1_b_bits_id; // @[Xbar.scala 231:30]
  wire [1:0] axi4xbar_auto_in_1_b_bits_resp; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_1_ar_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_1_ar_valid; // @[Xbar.scala 231:30]
  wire [5:0] axi4xbar_auto_in_1_ar_bits_id; // @[Xbar.scala 231:30]
  wire [33:0] axi4xbar_auto_in_1_ar_bits_addr; // @[Xbar.scala 231:30]
  wire [7:0] axi4xbar_auto_in_1_ar_bits_len; // @[Xbar.scala 231:30]
  wire [2:0] axi4xbar_auto_in_1_ar_bits_size; // @[Xbar.scala 231:30]
  wire [1:0] axi4xbar_auto_in_1_ar_bits_burst; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_1_ar_bits_lock; // @[Xbar.scala 231:30]
  wire [3:0] axi4xbar_auto_in_1_ar_bits_cache; // @[Xbar.scala 231:30]
  wire [2:0] axi4xbar_auto_in_1_ar_bits_prot; // @[Xbar.scala 231:30]
  wire [3:0] axi4xbar_auto_in_1_ar_bits_qos; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_1_r_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_1_r_valid; // @[Xbar.scala 231:30]
  wire [5:0] axi4xbar_auto_in_1_r_bits_id; // @[Xbar.scala 231:30]
  wire [511:0] axi4xbar_auto_in_1_r_bits_data; // @[Xbar.scala 231:30]
  wire [1:0] axi4xbar_auto_in_1_r_bits_resp; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_1_r_bits_last; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_0_aw_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_0_aw_valid; // @[Xbar.scala 231:30]
  wire [6:0] axi4xbar_auto_in_0_aw_bits_id; // @[Xbar.scala 231:30]
  wire [33:0] axi4xbar_auto_in_0_aw_bits_addr; // @[Xbar.scala 231:30]
  wire [7:0] axi4xbar_auto_in_0_aw_bits_len; // @[Xbar.scala 231:30]
  wire [2:0] axi4xbar_auto_in_0_aw_bits_size; // @[Xbar.scala 231:30]
  wire [1:0] axi4xbar_auto_in_0_aw_bits_burst; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_0_aw_bits_lock; // @[Xbar.scala 231:30]
  wire [3:0] axi4xbar_auto_in_0_aw_bits_cache; // @[Xbar.scala 231:30]
  wire [2:0] axi4xbar_auto_in_0_aw_bits_prot; // @[Xbar.scala 231:30]
  wire [3:0] axi4xbar_auto_in_0_aw_bits_qos; // @[Xbar.scala 231:30]
  wire [6:0] axi4xbar_auto_in_0_aw_bits_echo_tl_state_source; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_0_w_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_0_w_valid; // @[Xbar.scala 231:30]
  wire [511:0] axi4xbar_auto_in_0_w_bits_data; // @[Xbar.scala 231:30]
  wire [63:0] axi4xbar_auto_in_0_w_bits_strb; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_0_w_bits_last; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_0_b_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_0_b_valid; // @[Xbar.scala 231:30]
  wire [6:0] axi4xbar_auto_in_0_b_bits_id; // @[Xbar.scala 231:30]
  wire [6:0] axi4xbar_auto_in_0_b_bits_echo_tl_state_source; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_0_ar_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_0_ar_valid; // @[Xbar.scala 231:30]
  wire [6:0] axi4xbar_auto_in_0_ar_bits_id; // @[Xbar.scala 231:30]
  wire [33:0] axi4xbar_auto_in_0_ar_bits_addr; // @[Xbar.scala 231:30]
  wire [7:0] axi4xbar_auto_in_0_ar_bits_len; // @[Xbar.scala 231:30]
  wire [2:0] axi4xbar_auto_in_0_ar_bits_size; // @[Xbar.scala 231:30]
  wire [1:0] axi4xbar_auto_in_0_ar_bits_burst; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_0_ar_bits_lock; // @[Xbar.scala 231:30]
  wire [3:0] axi4xbar_auto_in_0_ar_bits_cache; // @[Xbar.scala 231:30]
  wire [2:0] axi4xbar_auto_in_0_ar_bits_prot; // @[Xbar.scala 231:30]
  wire [3:0] axi4xbar_auto_in_0_ar_bits_qos; // @[Xbar.scala 231:30]
  wire [6:0] axi4xbar_auto_in_0_ar_bits_echo_tl_state_source; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_0_r_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_0_r_valid; // @[Xbar.scala 231:30]
  wire [6:0] axi4xbar_auto_in_0_r_bits_id; // @[Xbar.scala 231:30]
  wire [511:0] axi4xbar_auto_in_0_r_bits_data; // @[Xbar.scala 231:30]
  wire [6:0] axi4xbar_auto_in_0_r_bits_echo_tl_state_source; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_in_0_r_bits_last; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_out_aw_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_out_aw_valid; // @[Xbar.scala 231:30]
  wire [7:0] axi4xbar_auto_out_aw_bits_id; // @[Xbar.scala 231:30]
  wire [33:0] axi4xbar_auto_out_aw_bits_addr; // @[Xbar.scala 231:30]
  wire [7:0] axi4xbar_auto_out_aw_bits_len; // @[Xbar.scala 231:30]
  wire [2:0] axi4xbar_auto_out_aw_bits_size; // @[Xbar.scala 231:30]
  wire [1:0] axi4xbar_auto_out_aw_bits_burst; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_out_aw_bits_lock; // @[Xbar.scala 231:30]
  wire [3:0] axi4xbar_auto_out_aw_bits_cache; // @[Xbar.scala 231:30]
  wire [2:0] axi4xbar_auto_out_aw_bits_prot; // @[Xbar.scala 231:30]
  wire [3:0] axi4xbar_auto_out_aw_bits_qos; // @[Xbar.scala 231:30]
  wire [6:0] axi4xbar_auto_out_aw_bits_echo_tl_state_source; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_out_w_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_out_w_valid; // @[Xbar.scala 231:30]
  wire [511:0] axi4xbar_auto_out_w_bits_data; // @[Xbar.scala 231:30]
  wire [63:0] axi4xbar_auto_out_w_bits_strb; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_out_w_bits_last; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_out_b_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_out_b_valid; // @[Xbar.scala 231:30]
  wire [7:0] axi4xbar_auto_out_b_bits_id; // @[Xbar.scala 231:30]
  wire [1:0] axi4xbar_auto_out_b_bits_resp; // @[Xbar.scala 231:30]
  wire [6:0] axi4xbar_auto_out_b_bits_echo_tl_state_source; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_out_ar_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_out_ar_valid; // @[Xbar.scala 231:30]
  wire [7:0] axi4xbar_auto_out_ar_bits_id; // @[Xbar.scala 231:30]
  wire [33:0] axi4xbar_auto_out_ar_bits_addr; // @[Xbar.scala 231:30]
  wire [7:0] axi4xbar_auto_out_ar_bits_len; // @[Xbar.scala 231:30]
  wire [2:0] axi4xbar_auto_out_ar_bits_size; // @[Xbar.scala 231:30]
  wire [1:0] axi4xbar_auto_out_ar_bits_burst; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_out_ar_bits_lock; // @[Xbar.scala 231:30]
  wire [3:0] axi4xbar_auto_out_ar_bits_cache; // @[Xbar.scala 231:30]
  wire [2:0] axi4xbar_auto_out_ar_bits_prot; // @[Xbar.scala 231:30]
  wire [3:0] axi4xbar_auto_out_ar_bits_qos; // @[Xbar.scala 231:30]
  wire [6:0] axi4xbar_auto_out_ar_bits_echo_tl_state_source; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_out_r_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_out_r_valid; // @[Xbar.scala 231:30]
  wire [7:0] axi4xbar_auto_out_r_bits_id; // @[Xbar.scala 231:30]
  wire [511:0] axi4xbar_auto_out_r_bits_data; // @[Xbar.scala 231:30]
  wire [1:0] axi4xbar_auto_out_r_bits_resp; // @[Xbar.scala 231:30]
  wire [6:0] axi4xbar_auto_out_r_bits_echo_tl_state_source; // @[Xbar.scala 231:30]
  wire  axi4xbar_auto_out_r_bits_last; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_clock; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_reset; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_in_aw_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_in_aw_valid; // @[Xbar.scala 231:30]
  wire [5:0] axi4xbar_1_auto_in_aw_bits_id; // @[Xbar.scala 231:30]
  wire [33:0] axi4xbar_1_auto_in_aw_bits_addr; // @[Xbar.scala 231:30]
  wire [7:0] axi4xbar_1_auto_in_aw_bits_len; // @[Xbar.scala 231:30]
  wire [2:0] axi4xbar_1_auto_in_aw_bits_size; // @[Xbar.scala 231:30]
  wire [1:0] axi4xbar_1_auto_in_aw_bits_burst; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_in_aw_bits_lock; // @[Xbar.scala 231:30]
  wire [3:0] axi4xbar_1_auto_in_aw_bits_cache; // @[Xbar.scala 231:30]
  wire [2:0] axi4xbar_1_auto_in_aw_bits_prot; // @[Xbar.scala 231:30]
  wire [3:0] axi4xbar_1_auto_in_aw_bits_qos; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_in_w_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_in_w_valid; // @[Xbar.scala 231:30]
  wire [511:0] axi4xbar_1_auto_in_w_bits_data; // @[Xbar.scala 231:30]
  wire [63:0] axi4xbar_1_auto_in_w_bits_strb; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_in_w_bits_last; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_in_b_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_in_b_valid; // @[Xbar.scala 231:30]
  wire [5:0] axi4xbar_1_auto_in_b_bits_id; // @[Xbar.scala 231:30]
  wire [1:0] axi4xbar_1_auto_in_b_bits_resp; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_in_ar_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_in_ar_valid; // @[Xbar.scala 231:30]
  wire [5:0] axi4xbar_1_auto_in_ar_bits_id; // @[Xbar.scala 231:30]
  wire [33:0] axi4xbar_1_auto_in_ar_bits_addr; // @[Xbar.scala 231:30]
  wire [7:0] axi4xbar_1_auto_in_ar_bits_len; // @[Xbar.scala 231:30]
  wire [2:0] axi4xbar_1_auto_in_ar_bits_size; // @[Xbar.scala 231:30]
  wire [1:0] axi4xbar_1_auto_in_ar_bits_burst; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_in_ar_bits_lock; // @[Xbar.scala 231:30]
  wire [3:0] axi4xbar_1_auto_in_ar_bits_cache; // @[Xbar.scala 231:30]
  wire [2:0] axi4xbar_1_auto_in_ar_bits_prot; // @[Xbar.scala 231:30]
  wire [3:0] axi4xbar_1_auto_in_ar_bits_qos; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_in_r_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_in_r_valid; // @[Xbar.scala 231:30]
  wire [5:0] axi4xbar_1_auto_in_r_bits_id; // @[Xbar.scala 231:30]
  wire [511:0] axi4xbar_1_auto_in_r_bits_data; // @[Xbar.scala 231:30]
  wire [1:0] axi4xbar_1_auto_in_r_bits_resp; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_in_r_bits_last; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_out_aw_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_out_aw_valid; // @[Xbar.scala 231:30]
  wire [5:0] axi4xbar_1_auto_out_aw_bits_id; // @[Xbar.scala 231:30]
  wire [33:0] axi4xbar_1_auto_out_aw_bits_addr; // @[Xbar.scala 231:30]
  wire [7:0] axi4xbar_1_auto_out_aw_bits_len; // @[Xbar.scala 231:30]
  wire [2:0] axi4xbar_1_auto_out_aw_bits_size; // @[Xbar.scala 231:30]
  wire [1:0] axi4xbar_1_auto_out_aw_bits_burst; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_out_aw_bits_lock; // @[Xbar.scala 231:30]
  wire [3:0] axi4xbar_1_auto_out_aw_bits_cache; // @[Xbar.scala 231:30]
  wire [2:0] axi4xbar_1_auto_out_aw_bits_prot; // @[Xbar.scala 231:30]
  wire [3:0] axi4xbar_1_auto_out_aw_bits_qos; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_out_w_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_out_w_valid; // @[Xbar.scala 231:30]
  wire [511:0] axi4xbar_1_auto_out_w_bits_data; // @[Xbar.scala 231:30]
  wire [63:0] axi4xbar_1_auto_out_w_bits_strb; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_out_w_bits_last; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_out_b_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_out_b_valid; // @[Xbar.scala 231:30]
  wire [5:0] axi4xbar_1_auto_out_b_bits_id; // @[Xbar.scala 231:30]
  wire [1:0] axi4xbar_1_auto_out_b_bits_resp; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_out_ar_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_out_ar_valid; // @[Xbar.scala 231:30]
  wire [5:0] axi4xbar_1_auto_out_ar_bits_id; // @[Xbar.scala 231:30]
  wire [33:0] axi4xbar_1_auto_out_ar_bits_addr; // @[Xbar.scala 231:30]
  wire [7:0] axi4xbar_1_auto_out_ar_bits_len; // @[Xbar.scala 231:30]
  wire [2:0] axi4xbar_1_auto_out_ar_bits_size; // @[Xbar.scala 231:30]
  wire [1:0] axi4xbar_1_auto_out_ar_bits_burst; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_out_ar_bits_lock; // @[Xbar.scala 231:30]
  wire [3:0] axi4xbar_1_auto_out_ar_bits_cache; // @[Xbar.scala 231:30]
  wire [2:0] axi4xbar_1_auto_out_ar_bits_prot; // @[Xbar.scala 231:30]
  wire [3:0] axi4xbar_1_auto_out_ar_bits_qos; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_out_r_ready; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_out_r_valid; // @[Xbar.scala 231:30]
  wire [5:0] axi4xbar_1_auto_out_r_bits_id; // @[Xbar.scala 231:30]
  wire [511:0] axi4xbar_1_auto_out_r_bits_data; // @[Xbar.scala 231:30]
  wire [1:0] axi4xbar_1_auto_out_r_bits_resp; // @[Xbar.scala 231:30]
  wire  axi4xbar_1_auto_out_r_bits_last; // @[Xbar.scala 231:30]
  wire  axi4buf_2_clock; // @[Buffer.scala 63:29]
  wire  axi4buf_2_reset; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_in_aw_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_in_aw_valid; // @[Buffer.scala 63:29]
  wire [5:0] axi4buf_2_auto_in_aw_bits_id; // @[Buffer.scala 63:29]
  wire [33:0] axi4buf_2_auto_in_aw_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_2_auto_in_aw_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_2_auto_in_aw_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_2_auto_in_aw_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_in_aw_bits_lock; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_2_auto_in_aw_bits_cache; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_2_auto_in_aw_bits_prot; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_2_auto_in_aw_bits_qos; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_in_w_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_in_w_valid; // @[Buffer.scala 63:29]
  wire [511:0] axi4buf_2_auto_in_w_bits_data; // @[Buffer.scala 63:29]
  wire [63:0] axi4buf_2_auto_in_w_bits_strb; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_in_w_bits_last; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_in_b_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_in_b_valid; // @[Buffer.scala 63:29]
  wire [5:0] axi4buf_2_auto_in_b_bits_id; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_2_auto_in_b_bits_resp; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_in_ar_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_in_ar_valid; // @[Buffer.scala 63:29]
  wire [5:0] axi4buf_2_auto_in_ar_bits_id; // @[Buffer.scala 63:29]
  wire [33:0] axi4buf_2_auto_in_ar_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_2_auto_in_ar_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_2_auto_in_ar_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_2_auto_in_ar_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_in_ar_bits_lock; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_2_auto_in_ar_bits_cache; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_2_auto_in_ar_bits_prot; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_2_auto_in_ar_bits_qos; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_in_r_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_in_r_valid; // @[Buffer.scala 63:29]
  wire [5:0] axi4buf_2_auto_in_r_bits_id; // @[Buffer.scala 63:29]
  wire [511:0] axi4buf_2_auto_in_r_bits_data; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_2_auto_in_r_bits_resp; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_in_r_bits_last; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_out_aw_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_out_aw_valid; // @[Buffer.scala 63:29]
  wire [5:0] axi4buf_2_auto_out_aw_bits_id; // @[Buffer.scala 63:29]
  wire [33:0] axi4buf_2_auto_out_aw_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_2_auto_out_aw_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_2_auto_out_aw_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_2_auto_out_aw_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_out_aw_bits_lock; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_2_auto_out_aw_bits_cache; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_2_auto_out_aw_bits_prot; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_2_auto_out_aw_bits_qos; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_out_w_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_out_w_valid; // @[Buffer.scala 63:29]
  wire [511:0] axi4buf_2_auto_out_w_bits_data; // @[Buffer.scala 63:29]
  wire [63:0] axi4buf_2_auto_out_w_bits_strb; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_out_w_bits_last; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_out_b_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_out_b_valid; // @[Buffer.scala 63:29]
  wire [5:0] axi4buf_2_auto_out_b_bits_id; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_2_auto_out_b_bits_resp; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_out_ar_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_out_ar_valid; // @[Buffer.scala 63:29]
  wire [5:0] axi4buf_2_auto_out_ar_bits_id; // @[Buffer.scala 63:29]
  wire [33:0] axi4buf_2_auto_out_ar_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_2_auto_out_ar_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_2_auto_out_ar_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_2_auto_out_ar_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_out_ar_bits_lock; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_2_auto_out_ar_bits_cache; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_2_auto_out_ar_bits_prot; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_2_auto_out_ar_bits_qos; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_out_r_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_out_r_valid; // @[Buffer.scala 63:29]
  wire [5:0] axi4buf_2_auto_out_r_bits_id; // @[Buffer.scala 63:29]
  wire [511:0] axi4buf_2_auto_out_r_bits_data; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_2_auto_out_r_bits_resp; // @[Buffer.scala 63:29]
  wire  axi4buf_2_auto_out_r_bits_last; // @[Buffer.scala 63:29]
  wire  axi4buf_3_clock; // @[Buffer.scala 63:29]
  wire  axi4buf_3_reset; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_in_aw_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_in_aw_valid; // @[Buffer.scala 63:29]
  wire [5:0] axi4buf_3_auto_in_aw_bits_id; // @[Buffer.scala 63:29]
  wire [33:0] axi4buf_3_auto_in_aw_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_3_auto_in_aw_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_3_auto_in_aw_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_3_auto_in_aw_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_in_aw_bits_lock; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_3_auto_in_aw_bits_cache; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_3_auto_in_aw_bits_prot; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_3_auto_in_aw_bits_qos; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_in_w_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_in_w_valid; // @[Buffer.scala 63:29]
  wire [511:0] axi4buf_3_auto_in_w_bits_data; // @[Buffer.scala 63:29]
  wire [63:0] axi4buf_3_auto_in_w_bits_strb; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_in_w_bits_last; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_in_b_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_in_b_valid; // @[Buffer.scala 63:29]
  wire [5:0] axi4buf_3_auto_in_b_bits_id; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_3_auto_in_b_bits_resp; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_in_ar_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_in_ar_valid; // @[Buffer.scala 63:29]
  wire [5:0] axi4buf_3_auto_in_ar_bits_id; // @[Buffer.scala 63:29]
  wire [33:0] axi4buf_3_auto_in_ar_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_3_auto_in_ar_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_3_auto_in_ar_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_3_auto_in_ar_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_in_ar_bits_lock; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_3_auto_in_ar_bits_cache; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_3_auto_in_ar_bits_prot; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_3_auto_in_ar_bits_qos; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_in_r_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_in_r_valid; // @[Buffer.scala 63:29]
  wire [5:0] axi4buf_3_auto_in_r_bits_id; // @[Buffer.scala 63:29]
  wire [511:0] axi4buf_3_auto_in_r_bits_data; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_3_auto_in_r_bits_resp; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_in_r_bits_last; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_out_aw_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_out_aw_valid; // @[Buffer.scala 63:29]
  wire [5:0] axi4buf_3_auto_out_aw_bits_id; // @[Buffer.scala 63:29]
  wire [33:0] axi4buf_3_auto_out_aw_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_3_auto_out_aw_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_3_auto_out_aw_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_3_auto_out_aw_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_out_aw_bits_lock; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_3_auto_out_aw_bits_cache; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_3_auto_out_aw_bits_prot; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_3_auto_out_aw_bits_qos; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_out_w_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_out_w_valid; // @[Buffer.scala 63:29]
  wire [511:0] axi4buf_3_auto_out_w_bits_data; // @[Buffer.scala 63:29]
  wire [63:0] axi4buf_3_auto_out_w_bits_strb; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_out_w_bits_last; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_out_b_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_out_b_valid; // @[Buffer.scala 63:29]
  wire [5:0] axi4buf_3_auto_out_b_bits_id; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_3_auto_out_b_bits_resp; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_out_ar_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_out_ar_valid; // @[Buffer.scala 63:29]
  wire [5:0] axi4buf_3_auto_out_ar_bits_id; // @[Buffer.scala 63:29]
  wire [33:0] axi4buf_3_auto_out_ar_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_3_auto_out_ar_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_3_auto_out_ar_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_3_auto_out_ar_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_out_ar_bits_lock; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_3_auto_out_ar_bits_cache; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_3_auto_out_ar_bits_prot; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_3_auto_out_ar_bits_qos; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_out_r_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_out_r_valid; // @[Buffer.scala 63:29]
  wire [5:0] axi4buf_3_auto_out_r_bits_id; // @[Buffer.scala 63:29]
  wire [511:0] axi4buf_3_auto_out_r_bits_data; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_3_auto_out_r_bits_resp; // @[Buffer.scala 63:29]
  wire  axi4buf_3_auto_out_r_bits_last; // @[Buffer.scala 63:29]
  wire  axi4yank_clock; // @[UserYanker.scala 108:30]
  wire  axi4yank_reset; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_aw_ready; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_aw_valid; // @[UserYanker.scala 108:30]
  wire [5:0] axi4yank_auto_in_aw_bits_id; // @[UserYanker.scala 108:30]
  wire [33:0] axi4yank_auto_in_aw_bits_addr; // @[UserYanker.scala 108:30]
  wire [7:0] axi4yank_auto_in_aw_bits_len; // @[UserYanker.scala 108:30]
  wire [2:0] axi4yank_auto_in_aw_bits_size; // @[UserYanker.scala 108:30]
  wire [1:0] axi4yank_auto_in_aw_bits_burst; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_aw_bits_lock; // @[UserYanker.scala 108:30]
  wire [3:0] axi4yank_auto_in_aw_bits_cache; // @[UserYanker.scala 108:30]
  wire [2:0] axi4yank_auto_in_aw_bits_prot; // @[UserYanker.scala 108:30]
  wire [3:0] axi4yank_auto_in_aw_bits_qos; // @[UserYanker.scala 108:30]
  wire [6:0] axi4yank_auto_in_aw_bits_echo_tl_state_source; // @[UserYanker.scala 108:30]
  wire [1:0] axi4yank_auto_in_aw_bits_echo_extra_id; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_w_ready; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_w_valid; // @[UserYanker.scala 108:30]
  wire [511:0] axi4yank_auto_in_w_bits_data; // @[UserYanker.scala 108:30]
  wire [63:0] axi4yank_auto_in_w_bits_strb; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_w_bits_last; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_b_ready; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_b_valid; // @[UserYanker.scala 108:30]
  wire [5:0] axi4yank_auto_in_b_bits_id; // @[UserYanker.scala 108:30]
  wire [1:0] axi4yank_auto_in_b_bits_resp; // @[UserYanker.scala 108:30]
  wire [6:0] axi4yank_auto_in_b_bits_echo_tl_state_source; // @[UserYanker.scala 108:30]
  wire [1:0] axi4yank_auto_in_b_bits_echo_extra_id; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_ar_ready; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_ar_valid; // @[UserYanker.scala 108:30]
  wire [5:0] axi4yank_auto_in_ar_bits_id; // @[UserYanker.scala 108:30]
  wire [33:0] axi4yank_auto_in_ar_bits_addr; // @[UserYanker.scala 108:30]
  wire [7:0] axi4yank_auto_in_ar_bits_len; // @[UserYanker.scala 108:30]
  wire [2:0] axi4yank_auto_in_ar_bits_size; // @[UserYanker.scala 108:30]
  wire [1:0] axi4yank_auto_in_ar_bits_burst; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_ar_bits_lock; // @[UserYanker.scala 108:30]
  wire [3:0] axi4yank_auto_in_ar_bits_cache; // @[UserYanker.scala 108:30]
  wire [2:0] axi4yank_auto_in_ar_bits_prot; // @[UserYanker.scala 108:30]
  wire [3:0] axi4yank_auto_in_ar_bits_qos; // @[UserYanker.scala 108:30]
  wire [6:0] axi4yank_auto_in_ar_bits_echo_tl_state_source; // @[UserYanker.scala 108:30]
  wire [1:0] axi4yank_auto_in_ar_bits_echo_extra_id; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_r_ready; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_r_valid; // @[UserYanker.scala 108:30]
  wire [5:0] axi4yank_auto_in_r_bits_id; // @[UserYanker.scala 108:30]
  wire [511:0] axi4yank_auto_in_r_bits_data; // @[UserYanker.scala 108:30]
  wire [1:0] axi4yank_auto_in_r_bits_resp; // @[UserYanker.scala 108:30]
  wire [6:0] axi4yank_auto_in_r_bits_echo_tl_state_source; // @[UserYanker.scala 108:30]
  wire [1:0] axi4yank_auto_in_r_bits_echo_extra_id; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_in_r_bits_last; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_aw_ready; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_aw_valid; // @[UserYanker.scala 108:30]
  wire [5:0] axi4yank_auto_out_aw_bits_id; // @[UserYanker.scala 108:30]
  wire [33:0] axi4yank_auto_out_aw_bits_addr; // @[UserYanker.scala 108:30]
  wire [7:0] axi4yank_auto_out_aw_bits_len; // @[UserYanker.scala 108:30]
  wire [2:0] axi4yank_auto_out_aw_bits_size; // @[UserYanker.scala 108:30]
  wire [1:0] axi4yank_auto_out_aw_bits_burst; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_aw_bits_lock; // @[UserYanker.scala 108:30]
  wire [3:0] axi4yank_auto_out_aw_bits_cache; // @[UserYanker.scala 108:30]
  wire [2:0] axi4yank_auto_out_aw_bits_prot; // @[UserYanker.scala 108:30]
  wire [3:0] axi4yank_auto_out_aw_bits_qos; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_w_ready; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_w_valid; // @[UserYanker.scala 108:30]
  wire [511:0] axi4yank_auto_out_w_bits_data; // @[UserYanker.scala 108:30]
  wire [63:0] axi4yank_auto_out_w_bits_strb; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_w_bits_last; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_b_ready; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_b_valid; // @[UserYanker.scala 108:30]
  wire [5:0] axi4yank_auto_out_b_bits_id; // @[UserYanker.scala 108:30]
  wire [1:0] axi4yank_auto_out_b_bits_resp; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_ar_ready; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_ar_valid; // @[UserYanker.scala 108:30]
  wire [5:0] axi4yank_auto_out_ar_bits_id; // @[UserYanker.scala 108:30]
  wire [33:0] axi4yank_auto_out_ar_bits_addr; // @[UserYanker.scala 108:30]
  wire [7:0] axi4yank_auto_out_ar_bits_len; // @[UserYanker.scala 108:30]
  wire [2:0] axi4yank_auto_out_ar_bits_size; // @[UserYanker.scala 108:30]
  wire [1:0] axi4yank_auto_out_ar_bits_burst; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_ar_bits_lock; // @[UserYanker.scala 108:30]
  wire [3:0] axi4yank_auto_out_ar_bits_cache; // @[UserYanker.scala 108:30]
  wire [2:0] axi4yank_auto_out_ar_bits_prot; // @[UserYanker.scala 108:30]
  wire [3:0] axi4yank_auto_out_ar_bits_qos; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_r_ready; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_r_valid; // @[UserYanker.scala 108:30]
  wire [5:0] axi4yank_auto_out_r_bits_id; // @[UserYanker.scala 108:30]
  wire [511:0] axi4yank_auto_out_r_bits_data; // @[UserYanker.scala 108:30]
  wire [1:0] axi4yank_auto_out_r_bits_resp; // @[UserYanker.scala 108:30]
  wire  axi4yank_auto_out_r_bits_last; // @[UserYanker.scala 108:30]
  wire  axi4buf_4_clock; // @[Buffer.scala 63:29]
  wire  axi4buf_4_reset; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_in_aw_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_in_aw_valid; // @[Buffer.scala 63:29]
  wire [5:0] axi4buf_4_auto_in_aw_bits_id; // @[Buffer.scala 63:29]
  wire [33:0] axi4buf_4_auto_in_aw_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_4_auto_in_aw_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_4_auto_in_aw_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_4_auto_in_aw_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_in_aw_bits_lock; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_4_auto_in_aw_bits_cache; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_4_auto_in_aw_bits_prot; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_4_auto_in_aw_bits_qos; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_4_auto_in_aw_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_4_auto_in_aw_bits_echo_extra_id; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_in_w_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_in_w_valid; // @[Buffer.scala 63:29]
  wire [511:0] axi4buf_4_auto_in_w_bits_data; // @[Buffer.scala 63:29]
  wire [63:0] axi4buf_4_auto_in_w_bits_strb; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_in_w_bits_last; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_in_b_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_in_b_valid; // @[Buffer.scala 63:29]
  wire [5:0] axi4buf_4_auto_in_b_bits_id; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_4_auto_in_b_bits_resp; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_4_auto_in_b_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_4_auto_in_b_bits_echo_extra_id; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_in_ar_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_in_ar_valid; // @[Buffer.scala 63:29]
  wire [5:0] axi4buf_4_auto_in_ar_bits_id; // @[Buffer.scala 63:29]
  wire [33:0] axi4buf_4_auto_in_ar_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_4_auto_in_ar_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_4_auto_in_ar_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_4_auto_in_ar_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_in_ar_bits_lock; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_4_auto_in_ar_bits_cache; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_4_auto_in_ar_bits_prot; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_4_auto_in_ar_bits_qos; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_4_auto_in_ar_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_4_auto_in_ar_bits_echo_extra_id; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_in_r_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_in_r_valid; // @[Buffer.scala 63:29]
  wire [5:0] axi4buf_4_auto_in_r_bits_id; // @[Buffer.scala 63:29]
  wire [511:0] axi4buf_4_auto_in_r_bits_data; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_4_auto_in_r_bits_resp; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_4_auto_in_r_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_4_auto_in_r_bits_echo_extra_id; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_in_r_bits_last; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_out_aw_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_out_aw_valid; // @[Buffer.scala 63:29]
  wire [5:0] axi4buf_4_auto_out_aw_bits_id; // @[Buffer.scala 63:29]
  wire [33:0] axi4buf_4_auto_out_aw_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_4_auto_out_aw_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_4_auto_out_aw_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_4_auto_out_aw_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_out_aw_bits_lock; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_4_auto_out_aw_bits_cache; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_4_auto_out_aw_bits_prot; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_4_auto_out_aw_bits_qos; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_4_auto_out_aw_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_4_auto_out_aw_bits_echo_extra_id; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_out_w_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_out_w_valid; // @[Buffer.scala 63:29]
  wire [511:0] axi4buf_4_auto_out_w_bits_data; // @[Buffer.scala 63:29]
  wire [63:0] axi4buf_4_auto_out_w_bits_strb; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_out_w_bits_last; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_out_b_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_out_b_valid; // @[Buffer.scala 63:29]
  wire [5:0] axi4buf_4_auto_out_b_bits_id; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_4_auto_out_b_bits_resp; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_4_auto_out_b_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_4_auto_out_b_bits_echo_extra_id; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_out_ar_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_out_ar_valid; // @[Buffer.scala 63:29]
  wire [5:0] axi4buf_4_auto_out_ar_bits_id; // @[Buffer.scala 63:29]
  wire [33:0] axi4buf_4_auto_out_ar_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_4_auto_out_ar_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_4_auto_out_ar_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_4_auto_out_ar_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_out_ar_bits_lock; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_4_auto_out_ar_bits_cache; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_4_auto_out_ar_bits_prot; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_4_auto_out_ar_bits_qos; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_4_auto_out_ar_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_4_auto_out_ar_bits_echo_extra_id; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_out_r_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_out_r_valid; // @[Buffer.scala 63:29]
  wire [5:0] axi4buf_4_auto_out_r_bits_id; // @[Buffer.scala 63:29]
  wire [511:0] axi4buf_4_auto_out_r_bits_data; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_4_auto_out_r_bits_resp; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_4_auto_out_r_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_4_auto_out_r_bits_echo_extra_id; // @[Buffer.scala 63:29]
  wire  axi4buf_4_auto_out_r_bits_last; // @[Buffer.scala 63:29]
  wire  axi4index_auto_in_aw_ready; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_in_aw_valid; // @[IdIndexer.scala 94:31]
  wire [7:0] axi4index_auto_in_aw_bits_id; // @[IdIndexer.scala 94:31]
  wire [33:0] axi4index_auto_in_aw_bits_addr; // @[IdIndexer.scala 94:31]
  wire [7:0] axi4index_auto_in_aw_bits_len; // @[IdIndexer.scala 94:31]
  wire [2:0] axi4index_auto_in_aw_bits_size; // @[IdIndexer.scala 94:31]
  wire [1:0] axi4index_auto_in_aw_bits_burst; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_in_aw_bits_lock; // @[IdIndexer.scala 94:31]
  wire [3:0] axi4index_auto_in_aw_bits_cache; // @[IdIndexer.scala 94:31]
  wire [2:0] axi4index_auto_in_aw_bits_prot; // @[IdIndexer.scala 94:31]
  wire [3:0] axi4index_auto_in_aw_bits_qos; // @[IdIndexer.scala 94:31]
  wire [6:0] axi4index_auto_in_aw_bits_echo_tl_state_source; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_in_w_ready; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_in_w_valid; // @[IdIndexer.scala 94:31]
  wire [511:0] axi4index_auto_in_w_bits_data; // @[IdIndexer.scala 94:31]
  wire [63:0] axi4index_auto_in_w_bits_strb; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_in_w_bits_last; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_in_b_ready; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_in_b_valid; // @[IdIndexer.scala 94:31]
  wire [7:0] axi4index_auto_in_b_bits_id; // @[IdIndexer.scala 94:31]
  wire [1:0] axi4index_auto_in_b_bits_resp; // @[IdIndexer.scala 94:31]
  wire [6:0] axi4index_auto_in_b_bits_echo_tl_state_source; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_in_ar_ready; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_in_ar_valid; // @[IdIndexer.scala 94:31]
  wire [7:0] axi4index_auto_in_ar_bits_id; // @[IdIndexer.scala 94:31]
  wire [33:0] axi4index_auto_in_ar_bits_addr; // @[IdIndexer.scala 94:31]
  wire [7:0] axi4index_auto_in_ar_bits_len; // @[IdIndexer.scala 94:31]
  wire [2:0] axi4index_auto_in_ar_bits_size; // @[IdIndexer.scala 94:31]
  wire [1:0] axi4index_auto_in_ar_bits_burst; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_in_ar_bits_lock; // @[IdIndexer.scala 94:31]
  wire [3:0] axi4index_auto_in_ar_bits_cache; // @[IdIndexer.scala 94:31]
  wire [2:0] axi4index_auto_in_ar_bits_prot; // @[IdIndexer.scala 94:31]
  wire [3:0] axi4index_auto_in_ar_bits_qos; // @[IdIndexer.scala 94:31]
  wire [6:0] axi4index_auto_in_ar_bits_echo_tl_state_source; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_in_r_ready; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_in_r_valid; // @[IdIndexer.scala 94:31]
  wire [7:0] axi4index_auto_in_r_bits_id; // @[IdIndexer.scala 94:31]
  wire [511:0] axi4index_auto_in_r_bits_data; // @[IdIndexer.scala 94:31]
  wire [1:0] axi4index_auto_in_r_bits_resp; // @[IdIndexer.scala 94:31]
  wire [6:0] axi4index_auto_in_r_bits_echo_tl_state_source; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_in_r_bits_last; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_aw_ready; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_aw_valid; // @[IdIndexer.scala 94:31]
  wire [5:0] axi4index_auto_out_aw_bits_id; // @[IdIndexer.scala 94:31]
  wire [33:0] axi4index_auto_out_aw_bits_addr; // @[IdIndexer.scala 94:31]
  wire [7:0] axi4index_auto_out_aw_bits_len; // @[IdIndexer.scala 94:31]
  wire [2:0] axi4index_auto_out_aw_bits_size; // @[IdIndexer.scala 94:31]
  wire [1:0] axi4index_auto_out_aw_bits_burst; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_aw_bits_lock; // @[IdIndexer.scala 94:31]
  wire [3:0] axi4index_auto_out_aw_bits_cache; // @[IdIndexer.scala 94:31]
  wire [2:0] axi4index_auto_out_aw_bits_prot; // @[IdIndexer.scala 94:31]
  wire [3:0] axi4index_auto_out_aw_bits_qos; // @[IdIndexer.scala 94:31]
  wire [6:0] axi4index_auto_out_aw_bits_echo_tl_state_source; // @[IdIndexer.scala 94:31]
  wire [1:0] axi4index_auto_out_aw_bits_echo_extra_id; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_w_ready; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_w_valid; // @[IdIndexer.scala 94:31]
  wire [511:0] axi4index_auto_out_w_bits_data; // @[IdIndexer.scala 94:31]
  wire [63:0] axi4index_auto_out_w_bits_strb; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_w_bits_last; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_b_ready; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_b_valid; // @[IdIndexer.scala 94:31]
  wire [5:0] axi4index_auto_out_b_bits_id; // @[IdIndexer.scala 94:31]
  wire [1:0] axi4index_auto_out_b_bits_resp; // @[IdIndexer.scala 94:31]
  wire [6:0] axi4index_auto_out_b_bits_echo_tl_state_source; // @[IdIndexer.scala 94:31]
  wire [1:0] axi4index_auto_out_b_bits_echo_extra_id; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_ar_ready; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_ar_valid; // @[IdIndexer.scala 94:31]
  wire [5:0] axi4index_auto_out_ar_bits_id; // @[IdIndexer.scala 94:31]
  wire [33:0] axi4index_auto_out_ar_bits_addr; // @[IdIndexer.scala 94:31]
  wire [7:0] axi4index_auto_out_ar_bits_len; // @[IdIndexer.scala 94:31]
  wire [2:0] axi4index_auto_out_ar_bits_size; // @[IdIndexer.scala 94:31]
  wire [1:0] axi4index_auto_out_ar_bits_burst; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_ar_bits_lock; // @[IdIndexer.scala 94:31]
  wire [3:0] axi4index_auto_out_ar_bits_cache; // @[IdIndexer.scala 94:31]
  wire [2:0] axi4index_auto_out_ar_bits_prot; // @[IdIndexer.scala 94:31]
  wire [3:0] axi4index_auto_out_ar_bits_qos; // @[IdIndexer.scala 94:31]
  wire [6:0] axi4index_auto_out_ar_bits_echo_tl_state_source; // @[IdIndexer.scala 94:31]
  wire [1:0] axi4index_auto_out_ar_bits_echo_extra_id; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_r_ready; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_r_valid; // @[IdIndexer.scala 94:31]
  wire [5:0] axi4index_auto_out_r_bits_id; // @[IdIndexer.scala 94:31]
  wire [511:0] axi4index_auto_out_r_bits_data; // @[IdIndexer.scala 94:31]
  wire [1:0] axi4index_auto_out_r_bits_resp; // @[IdIndexer.scala 94:31]
  wire [6:0] axi4index_auto_out_r_bits_echo_tl_state_source; // @[IdIndexer.scala 94:31]
  wire [1:0] axi4index_auto_out_r_bits_echo_extra_id; // @[IdIndexer.scala 94:31]
  wire  axi4index_auto_out_r_bits_last; // @[IdIndexer.scala 94:31]
  wire  axi4buf_5_clock; // @[Buffer.scala 63:29]
  wire  axi4buf_5_reset; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_in_aw_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_in_aw_valid; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_5_auto_in_aw_bits_id; // @[Buffer.scala 63:29]
  wire [33:0] axi4buf_5_auto_in_aw_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_5_auto_in_aw_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_5_auto_in_aw_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_5_auto_in_aw_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_in_aw_bits_lock; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_5_auto_in_aw_bits_cache; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_5_auto_in_aw_bits_prot; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_5_auto_in_aw_bits_qos; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_5_auto_in_aw_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_in_w_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_in_w_valid; // @[Buffer.scala 63:29]
  wire [511:0] axi4buf_5_auto_in_w_bits_data; // @[Buffer.scala 63:29]
  wire [63:0] axi4buf_5_auto_in_w_bits_strb; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_in_w_bits_last; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_in_b_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_in_b_valid; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_5_auto_in_b_bits_id; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_5_auto_in_b_bits_resp; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_5_auto_in_b_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_in_ar_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_in_ar_valid; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_5_auto_in_ar_bits_id; // @[Buffer.scala 63:29]
  wire [33:0] axi4buf_5_auto_in_ar_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_5_auto_in_ar_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_5_auto_in_ar_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_5_auto_in_ar_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_in_ar_bits_lock; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_5_auto_in_ar_bits_cache; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_5_auto_in_ar_bits_prot; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_5_auto_in_ar_bits_qos; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_5_auto_in_ar_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_in_r_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_in_r_valid; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_5_auto_in_r_bits_id; // @[Buffer.scala 63:29]
  wire [511:0] axi4buf_5_auto_in_r_bits_data; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_5_auto_in_r_bits_resp; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_5_auto_in_r_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_in_r_bits_last; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_out_aw_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_out_aw_valid; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_5_auto_out_aw_bits_id; // @[Buffer.scala 63:29]
  wire [33:0] axi4buf_5_auto_out_aw_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_5_auto_out_aw_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_5_auto_out_aw_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_5_auto_out_aw_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_out_aw_bits_lock; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_5_auto_out_aw_bits_cache; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_5_auto_out_aw_bits_prot; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_5_auto_out_aw_bits_qos; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_5_auto_out_aw_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_out_w_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_out_w_valid; // @[Buffer.scala 63:29]
  wire [511:0] axi4buf_5_auto_out_w_bits_data; // @[Buffer.scala 63:29]
  wire [63:0] axi4buf_5_auto_out_w_bits_strb; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_out_w_bits_last; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_out_b_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_out_b_valid; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_5_auto_out_b_bits_id; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_5_auto_out_b_bits_resp; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_5_auto_out_b_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_out_ar_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_out_ar_valid; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_5_auto_out_ar_bits_id; // @[Buffer.scala 63:29]
  wire [33:0] axi4buf_5_auto_out_ar_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_5_auto_out_ar_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_5_auto_out_ar_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_5_auto_out_ar_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_out_ar_bits_lock; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_5_auto_out_ar_bits_cache; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_5_auto_out_ar_bits_prot; // @[Buffer.scala 63:29]
  wire [3:0] axi4buf_5_auto_out_ar_bits_qos; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_5_auto_out_ar_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_out_r_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_out_r_valid; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_5_auto_out_r_bits_id; // @[Buffer.scala 63:29]
  wire [511:0] axi4buf_5_auto_out_r_bits_data; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_5_auto_out_r_bits_resp; // @[Buffer.scala 63:29]
  wire [6:0] axi4buf_5_auto_out_r_bits_echo_tl_state_source; // @[Buffer.scala 63:29]
  wire  axi4buf_5_auto_out_r_bits_last; // @[Buffer.scala 63:29]
  wire  cmd_resp_axilhub_clock; // @[ComposerTop.scala 134:36]
  wire  cmd_resp_axilhub_reset; // @[ComposerTop.scala 134:36]
  wire  cmd_resp_axilhub_auto_in_aw_ready; // @[ComposerTop.scala 134:36]
  wire  cmd_resp_axilhub_auto_in_aw_valid; // @[ComposerTop.scala 134:36]
  wire [15:0] cmd_resp_axilhub_auto_in_aw_bits_id; // @[ComposerTop.scala 134:36]
  wire [15:0] cmd_resp_axilhub_auto_in_aw_bits_addr; // @[ComposerTop.scala 134:36]
  wire [7:0] cmd_resp_axilhub_auto_in_aw_bits_len; // @[ComposerTop.scala 134:36]
  wire [2:0] cmd_resp_axilhub_auto_in_aw_bits_size; // @[ComposerTop.scala 134:36]
  wire [1:0] cmd_resp_axilhub_auto_in_aw_bits_burst; // @[ComposerTop.scala 134:36]
  wire  cmd_resp_axilhub_auto_in_w_ready; // @[ComposerTop.scala 134:36]
  wire  cmd_resp_axilhub_auto_in_w_valid; // @[ComposerTop.scala 134:36]
  wire [31:0] cmd_resp_axilhub_auto_in_w_bits_data; // @[ComposerTop.scala 134:36]
  wire  cmd_resp_axilhub_auto_in_w_bits_last; // @[ComposerTop.scala 134:36]
  wire  cmd_resp_axilhub_auto_in_b_ready; // @[ComposerTop.scala 134:36]
  wire  cmd_resp_axilhub_auto_in_b_valid; // @[ComposerTop.scala 134:36]
  wire [15:0] cmd_resp_axilhub_auto_in_b_bits_id; // @[ComposerTop.scala 134:36]
  wire [1:0] cmd_resp_axilhub_auto_in_b_bits_resp; // @[ComposerTop.scala 134:36]
  wire  cmd_resp_axilhub_auto_in_ar_ready; // @[ComposerTop.scala 134:36]
  wire  cmd_resp_axilhub_auto_in_ar_valid; // @[ComposerTop.scala 134:36]
  wire [15:0] cmd_resp_axilhub_auto_in_ar_bits_id; // @[ComposerTop.scala 134:36]
  wire [15:0] cmd_resp_axilhub_auto_in_ar_bits_addr; // @[ComposerTop.scala 134:36]
  wire [7:0] cmd_resp_axilhub_auto_in_ar_bits_len; // @[ComposerTop.scala 134:36]
  wire [2:0] cmd_resp_axilhub_auto_in_ar_bits_size; // @[ComposerTop.scala 134:36]
  wire [1:0] cmd_resp_axilhub_auto_in_ar_bits_burst; // @[ComposerTop.scala 134:36]
  wire  cmd_resp_axilhub_auto_in_r_ready; // @[ComposerTop.scala 134:36]
  wire  cmd_resp_axilhub_auto_in_r_valid; // @[ComposerTop.scala 134:36]
  wire [15:0] cmd_resp_axilhub_auto_in_r_bits_id; // @[ComposerTop.scala 134:36]
  wire [31:0] cmd_resp_axilhub_auto_in_r_bits_data; // @[ComposerTop.scala 134:36]
  wire [1:0] cmd_resp_axilhub_auto_in_r_bits_resp; // @[ComposerTop.scala 134:36]
  wire  cmd_resp_axilhub_auto_in_r_bits_last; // @[ComposerTop.scala 134:36]
  wire  cmd_resp_axilhub_io_rocc_in_ready; // @[ComposerTop.scala 134:36]
  wire  cmd_resp_axilhub_io_rocc_in_valid; // @[ComposerTop.scala 134:36]
  wire [6:0] cmd_resp_axilhub_io_rocc_in_bits_inst_funct; // @[ComposerTop.scala 134:36]
  wire [4:0] cmd_resp_axilhub_io_rocc_in_bits_inst_rs2; // @[ComposerTop.scala 134:36]
  wire [4:0] cmd_resp_axilhub_io_rocc_in_bits_inst_rs1; // @[ComposerTop.scala 134:36]
  wire [6:0] cmd_resp_axilhub_io_rocc_in_bits_inst_opcode; // @[ComposerTop.scala 134:36]
  wire [63:0] cmd_resp_axilhub_io_rocc_in_bits_rs1; // @[ComposerTop.scala 134:36]
  wire [63:0] cmd_resp_axilhub_io_rocc_in_bits_rs2; // @[ComposerTop.scala 134:36]
  wire  cmd_resp_axilhub_io_rocc_out_ready; // @[ComposerTop.scala 134:36]
  wire  cmd_resp_axilhub_io_rocc_out_valid; // @[ComposerTop.scala 134:36]
  wire [4:0] cmd_resp_axilhub_io_rocc_out_bits_rd; // @[ComposerTop.scala 134:36]
  wire [63:0] cmd_resp_axilhub_io_rocc_out_bits_data; // @[ComposerTop.scala 134:36]
  wire  axi4buf_6_clock; // @[Buffer.scala 63:29]
  wire  axi4buf_6_reset; // @[Buffer.scala 63:29]
  wire  axi4buf_6_auto_in_aw_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_6_auto_in_aw_valid; // @[Buffer.scala 63:29]
  wire [15:0] axi4buf_6_auto_in_aw_bits_id; // @[Buffer.scala 63:29]
  wire [15:0] axi4buf_6_auto_in_aw_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_6_auto_in_aw_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_6_auto_in_aw_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_6_auto_in_aw_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_6_auto_in_w_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_6_auto_in_w_valid; // @[Buffer.scala 63:29]
  wire [31:0] axi4buf_6_auto_in_w_bits_data; // @[Buffer.scala 63:29]
  wire  axi4buf_6_auto_in_w_bits_last; // @[Buffer.scala 63:29]
  wire  axi4buf_6_auto_in_b_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_6_auto_in_b_valid; // @[Buffer.scala 63:29]
  wire [15:0] axi4buf_6_auto_in_b_bits_id; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_6_auto_in_b_bits_resp; // @[Buffer.scala 63:29]
  wire  axi4buf_6_auto_in_ar_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_6_auto_in_ar_valid; // @[Buffer.scala 63:29]
  wire [15:0] axi4buf_6_auto_in_ar_bits_id; // @[Buffer.scala 63:29]
  wire [15:0] axi4buf_6_auto_in_ar_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_6_auto_in_ar_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_6_auto_in_ar_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_6_auto_in_ar_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_6_auto_in_r_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_6_auto_in_r_valid; // @[Buffer.scala 63:29]
  wire [15:0] axi4buf_6_auto_in_r_bits_id; // @[Buffer.scala 63:29]
  wire [31:0] axi4buf_6_auto_in_r_bits_data; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_6_auto_in_r_bits_resp; // @[Buffer.scala 63:29]
  wire  axi4buf_6_auto_in_r_bits_last; // @[Buffer.scala 63:29]
  wire  axi4buf_6_auto_out_aw_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_6_auto_out_aw_valid; // @[Buffer.scala 63:29]
  wire [15:0] axi4buf_6_auto_out_aw_bits_id; // @[Buffer.scala 63:29]
  wire [15:0] axi4buf_6_auto_out_aw_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_6_auto_out_aw_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_6_auto_out_aw_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_6_auto_out_aw_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_6_auto_out_w_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_6_auto_out_w_valid; // @[Buffer.scala 63:29]
  wire [31:0] axi4buf_6_auto_out_w_bits_data; // @[Buffer.scala 63:29]
  wire  axi4buf_6_auto_out_w_bits_last; // @[Buffer.scala 63:29]
  wire  axi4buf_6_auto_out_b_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_6_auto_out_b_valid; // @[Buffer.scala 63:29]
  wire [15:0] axi4buf_6_auto_out_b_bits_id; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_6_auto_out_b_bits_resp; // @[Buffer.scala 63:29]
  wire  axi4buf_6_auto_out_ar_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_6_auto_out_ar_valid; // @[Buffer.scala 63:29]
  wire [15:0] axi4buf_6_auto_out_ar_bits_id; // @[Buffer.scala 63:29]
  wire [15:0] axi4buf_6_auto_out_ar_bits_addr; // @[Buffer.scala 63:29]
  wire [7:0] axi4buf_6_auto_out_ar_bits_len; // @[Buffer.scala 63:29]
  wire [2:0] axi4buf_6_auto_out_ar_bits_size; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_6_auto_out_ar_bits_burst; // @[Buffer.scala 63:29]
  wire  axi4buf_6_auto_out_r_ready; // @[Buffer.scala 63:29]
  wire  axi4buf_6_auto_out_r_valid; // @[Buffer.scala 63:29]
  wire [15:0] axi4buf_6_auto_out_r_bits_id; // @[Buffer.scala 63:29]
  wire [31:0] axi4buf_6_auto_out_r_bits_data; // @[Buffer.scala 63:29]
  wire [1:0] axi4buf_6_auto_out_r_bits_resp; // @[Buffer.scala 63:29]
  wire  axi4buf_6_auto_out_r_bits_last; // @[Buffer.scala 63:29]
  reg [63:0] arCnt; // @[ComposerTop.scala 171:22]
  reg [63:0] awCnt; // @[ComposerTop.scala 172:22]
  reg [63:0] rCnt; // @[ComposerTop.scala 173:21]
  reg [63:0] wCnt; // @[ComposerTop.scala 174:21]
  reg [63:0] bCnt; // @[ComposerTop.scala 175:21]
  wire  q_ar_valid = axi4buf_3_auto_out_ar_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire  _T = M00_AXI_arready & q_ar_valid; // @[Decoupled.scala 51:35]
  wire [63:0] _arCnt_T_1 = arCnt + 64'h1; // @[ComposerTop.scala 179:20]
  wire  q_aw_valid = axi4buf_3_auto_out_aw_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire  _T_1 = M00_AXI_awready & q_aw_valid; // @[Decoupled.scala 51:35]
  wire [63:0] _awCnt_T_1 = awCnt + 64'h1; // @[ComposerTop.scala 182:20]
  wire  q_r_ready = axi4buf_3_auto_out_r_ready; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire  _T_2 = q_r_ready & M00_AXI_rvalid; // @[Decoupled.scala 51:35]
  wire [63:0] _rCnt_T_1 = rCnt + 64'h1; // @[ComposerTop.scala 185:18]
  wire  q_w_valid = axi4buf_3_auto_out_w_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire  _T_3 = M00_AXI_wready & q_w_valid; // @[Decoupled.scala 51:35]
  wire [63:0] _wCnt_T_1 = wCnt + 64'h1; // @[ComposerTop.scala 188:18]
  wire  q_b_ready = axi4buf_3_auto_out_b_ready; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire  _T_4 = q_b_ready & M00_AXI_bvalid; // @[Decoupled.scala 51:35]
  wire [63:0] _bCnt_T_1 = bCnt + 64'h1; // @[ComposerTop.scala 191:18]
  reg [63:0] rWait; // @[ComposerTop.scala 194:22]
  reg [63:0] bWait; // @[ComposerTop.scala 195:22]
  wire [63:0] _rWait_T_1 = rWait + 64'h1; // @[ComposerTop.scala 197:20]
  wire [63:0] _bWait_T_1 = bWait + 64'h1; // @[ComposerTop.scala 201:20]
  wire [63:0] _GEN_7 = 5'h16 == acc_io_resp_bits_rd ? bWait : acc_io_resp_bits_data; // @[ComposerTop.scala 149:31 204:38 224:45]
  wire [63:0] _GEN_8 = 5'h15 == acc_io_resp_bits_rd ? rWait : _GEN_7; // @[ComposerTop.scala 204:38 221:45]
  wire [63:0] _GEN_9 = 5'h14 == acc_io_resp_bits_rd ? bCnt : _GEN_8; // @[ComposerTop.scala 204:38 218:45]
  wire [63:0] _GEN_10 = 5'h13 == acc_io_resp_bits_rd ? wCnt : _GEN_9; // @[ComposerTop.scala 204:38 215:45]
  wire [63:0] _GEN_11 = 5'h12 == acc_io_resp_bits_rd ? rCnt : _GEN_10; // @[ComposerTop.scala 204:38 212:45]
  wire [63:0] _GEN_12 = 5'h11 == acc_io_resp_bits_rd ? awCnt : _GEN_11; // @[ComposerTop.scala 204:38 209:45]
  ComposerAccSystem acc ( // @[ComposerTop.scala 80:23]
    .clock(acc_clock),
    .reset(acc_reset),
    .auto_mem_out_a_ready(acc_auto_mem_out_a_ready),
    .auto_mem_out_a_valid(acc_auto_mem_out_a_valid),
    .auto_mem_out_a_bits_opcode(acc_auto_mem_out_a_bits_opcode),
    .auto_mem_out_a_bits_size(acc_auto_mem_out_a_bits_size),
    .auto_mem_out_a_bits_source(acc_auto_mem_out_a_bits_source),
    .auto_mem_out_a_bits_address(acc_auto_mem_out_a_bits_address),
    .auto_mem_out_a_bits_mask(acc_auto_mem_out_a_bits_mask),
    .auto_mem_out_a_bits_data(acc_auto_mem_out_a_bits_data),
    .auto_mem_out_d_ready(acc_auto_mem_out_d_ready),
    .auto_mem_out_d_valid(acc_auto_mem_out_d_valid),
    .auto_mem_out_d_bits_source(acc_auto_mem_out_d_bits_source),
    .auto_mem_out_d_bits_data(acc_auto_mem_out_d_bits_data),
    .io_cmd_ready(acc_io_cmd_ready),
    .io_cmd_valid(acc_io_cmd_valid),
    .io_cmd_bits_inst_funct(acc_io_cmd_bits_inst_funct),
    .io_cmd_bits_inst_rs2(acc_io_cmd_bits_inst_rs2),
    .io_cmd_bits_inst_rs1(acc_io_cmd_bits_inst_rs1),
    .io_cmd_bits_inst_opcode(acc_io_cmd_bits_inst_opcode),
    .io_cmd_bits_rs1(acc_io_cmd_bits_rs1),
    .io_cmd_bits_rs2(acc_io_cmd_bits_rs2),
    .io_resp_ready(acc_io_resp_ready),
    .io_resp_valid(acc_io_resp_valid),
    .io_resp_bits_rd(acc_io_resp_bits_rd),
    .io_resp_bits_data(acc_io_resp_bits_data)
  );
  AXI4Buffer axi4buf ( // @[Buffer.scala 63:29]
    .clock(axi4buf_clock),
    .reset(axi4buf_reset),
    .auto_in_aw_ready(axi4buf_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4buf_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4buf_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axi4buf_auto_in_aw_bits_burst),
    .auto_in_aw_bits_lock(axi4buf_auto_in_aw_bits_lock),
    .auto_in_aw_bits_cache(axi4buf_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(axi4buf_auto_in_aw_bits_prot),
    .auto_in_aw_bits_qos(axi4buf_auto_in_aw_bits_qos),
    .auto_in_aw_bits_echo_tl_state_source(axi4buf_auto_in_aw_bits_echo_tl_state_source),
    .auto_in_w_ready(axi4buf_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_auto_in_b_bits_id),
    .auto_in_b_bits_echo_tl_state_source(axi4buf_auto_in_b_bits_echo_tl_state_source),
    .auto_in_ar_ready(axi4buf_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4buf_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4buf_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axi4buf_auto_in_ar_bits_burst),
    .auto_in_ar_bits_lock(axi4buf_auto_in_ar_bits_lock),
    .auto_in_ar_bits_cache(axi4buf_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(axi4buf_auto_in_ar_bits_prot),
    .auto_in_ar_bits_qos(axi4buf_auto_in_ar_bits_qos),
    .auto_in_ar_bits_echo_tl_state_source(axi4buf_auto_in_ar_bits_echo_tl_state_source),
    .auto_in_r_ready(axi4buf_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_auto_in_r_bits_data),
    .auto_in_r_bits_echo_tl_state_source(axi4buf_auto_in_r_bits_echo_tl_state_source),
    .auto_in_r_bits_last(axi4buf_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4buf_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4buf_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(axi4buf_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(axi4buf_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(axi4buf_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(axi4buf_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(axi4buf_auto_out_aw_bits_qos),
    .auto_out_aw_bits_echo_tl_state_source(axi4buf_auto_out_aw_bits_echo_tl_state_source),
    .auto_out_w_ready(axi4buf_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_auto_out_b_bits_id),
    .auto_out_b_bits_echo_tl_state_source(axi4buf_auto_out_b_bits_echo_tl_state_source),
    .auto_out_ar_ready(axi4buf_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4buf_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4buf_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(axi4buf_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(axi4buf_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(axi4buf_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(axi4buf_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(axi4buf_auto_out_ar_bits_qos),
    .auto_out_ar_bits_echo_tl_state_source(axi4buf_auto_out_ar_bits_echo_tl_state_source),
    .auto_out_r_ready(axi4buf_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_auto_out_r_bits_data),
    .auto_out_r_bits_echo_tl_state_source(axi4buf_auto_out_r_bits_echo_tl_state_source),
    .auto_out_r_bits_last(axi4buf_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_1 ( // @[Buffer.scala 63:29]
    .clock(axi4buf_1_clock),
    .reset(axi4buf_1_reset),
    .auto_in_aw_ready(axi4buf_1_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_1_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_1_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_1_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4buf_1_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4buf_1_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axi4buf_1_auto_in_aw_bits_burst),
    .auto_in_aw_bits_lock(axi4buf_1_auto_in_aw_bits_lock),
    .auto_in_aw_bits_cache(axi4buf_1_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(axi4buf_1_auto_in_aw_bits_prot),
    .auto_in_aw_bits_qos(axi4buf_1_auto_in_aw_bits_qos),
    .auto_in_aw_bits_echo_tl_state_source(axi4buf_1_auto_in_aw_bits_echo_tl_state_source),
    .auto_in_w_ready(axi4buf_1_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_1_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_1_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_1_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_1_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_1_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_1_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_1_auto_in_b_bits_id),
    .auto_in_b_bits_echo_tl_state_source(axi4buf_1_auto_in_b_bits_echo_tl_state_source),
    .auto_in_ar_ready(axi4buf_1_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_1_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_1_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_1_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4buf_1_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4buf_1_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axi4buf_1_auto_in_ar_bits_burst),
    .auto_in_ar_bits_lock(axi4buf_1_auto_in_ar_bits_lock),
    .auto_in_ar_bits_cache(axi4buf_1_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(axi4buf_1_auto_in_ar_bits_prot),
    .auto_in_ar_bits_qos(axi4buf_1_auto_in_ar_bits_qos),
    .auto_in_ar_bits_echo_tl_state_source(axi4buf_1_auto_in_ar_bits_echo_tl_state_source),
    .auto_in_r_ready(axi4buf_1_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_1_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_1_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_1_auto_in_r_bits_data),
    .auto_in_r_bits_echo_tl_state_source(axi4buf_1_auto_in_r_bits_echo_tl_state_source),
    .auto_in_r_bits_last(axi4buf_1_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_1_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_1_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_1_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_1_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4buf_1_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4buf_1_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(axi4buf_1_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(axi4buf_1_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(axi4buf_1_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(axi4buf_1_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(axi4buf_1_auto_out_aw_bits_qos),
    .auto_out_aw_bits_echo_tl_state_source(axi4buf_1_auto_out_aw_bits_echo_tl_state_source),
    .auto_out_w_ready(axi4buf_1_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_1_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_1_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_1_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_1_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_1_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_1_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_1_auto_out_b_bits_id),
    .auto_out_b_bits_echo_tl_state_source(axi4buf_1_auto_out_b_bits_echo_tl_state_source),
    .auto_out_ar_ready(axi4buf_1_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_1_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_1_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_1_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4buf_1_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4buf_1_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(axi4buf_1_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(axi4buf_1_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(axi4buf_1_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(axi4buf_1_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(axi4buf_1_auto_out_ar_bits_qos),
    .auto_out_ar_bits_echo_tl_state_source(axi4buf_1_auto_out_ar_bits_echo_tl_state_source),
    .auto_out_r_ready(axi4buf_1_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_1_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_1_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_1_auto_out_r_bits_data),
    .auto_out_r_bits_echo_tl_state_source(axi4buf_1_auto_out_r_bits_echo_tl_state_source),
    .auto_out_r_bits_last(axi4buf_1_auto_out_r_bits_last)
  );
  TLToAXI4 tl2axi4 ( // @[ToAXI4.scala 286:29]
    .clock(tl2axi4_clock),
    .reset(tl2axi4_reset),
    .auto_in_a_ready(tl2axi4_auto_in_a_ready),
    .auto_in_a_valid(tl2axi4_auto_in_a_valid),
    .auto_in_a_bits_opcode(tl2axi4_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(tl2axi4_auto_in_a_bits_size),
    .auto_in_a_bits_source(tl2axi4_auto_in_a_bits_source),
    .auto_in_a_bits_address(tl2axi4_auto_in_a_bits_address),
    .auto_in_a_bits_mask(tl2axi4_auto_in_a_bits_mask),
    .auto_in_a_bits_data(tl2axi4_auto_in_a_bits_data),
    .auto_in_d_ready(tl2axi4_auto_in_d_ready),
    .auto_in_d_valid(tl2axi4_auto_in_d_valid),
    .auto_in_d_bits_source(tl2axi4_auto_in_d_bits_source),
    .auto_in_d_bits_data(tl2axi4_auto_in_d_bits_data),
    .auto_out_aw_ready(tl2axi4_auto_out_aw_ready),
    .auto_out_aw_valid(tl2axi4_auto_out_aw_valid),
    .auto_out_aw_bits_id(tl2axi4_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(tl2axi4_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(tl2axi4_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(tl2axi4_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(tl2axi4_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(tl2axi4_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(tl2axi4_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(tl2axi4_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(tl2axi4_auto_out_aw_bits_qos),
    .auto_out_aw_bits_echo_tl_state_source(tl2axi4_auto_out_aw_bits_echo_tl_state_source),
    .auto_out_w_ready(tl2axi4_auto_out_w_ready),
    .auto_out_w_valid(tl2axi4_auto_out_w_valid),
    .auto_out_w_bits_data(tl2axi4_auto_out_w_bits_data),
    .auto_out_w_bits_strb(tl2axi4_auto_out_w_bits_strb),
    .auto_out_w_bits_last(tl2axi4_auto_out_w_bits_last),
    .auto_out_b_ready(tl2axi4_auto_out_b_ready),
    .auto_out_b_valid(tl2axi4_auto_out_b_valid),
    .auto_out_b_bits_id(tl2axi4_auto_out_b_bits_id),
    .auto_out_b_bits_echo_tl_state_source(tl2axi4_auto_out_b_bits_echo_tl_state_source),
    .auto_out_ar_ready(tl2axi4_auto_out_ar_ready),
    .auto_out_ar_valid(tl2axi4_auto_out_ar_valid),
    .auto_out_ar_bits_id(tl2axi4_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(tl2axi4_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(tl2axi4_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(tl2axi4_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(tl2axi4_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(tl2axi4_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(tl2axi4_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(tl2axi4_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(tl2axi4_auto_out_ar_bits_qos),
    .auto_out_ar_bits_echo_tl_state_source(tl2axi4_auto_out_ar_bits_echo_tl_state_source),
    .auto_out_r_ready(tl2axi4_auto_out_r_ready),
    .auto_out_r_valid(tl2axi4_auto_out_r_valid),
    .auto_out_r_bits_id(tl2axi4_auto_out_r_bits_id),
    .auto_out_r_bits_data(tl2axi4_auto_out_r_bits_data),
    .auto_out_r_bits_echo_tl_state_source(tl2axi4_auto_out_r_bits_echo_tl_state_source),
    .auto_out_r_bits_last(tl2axi4_auto_out_r_bits_last)
  );
  AXI4Xbar axi4xbar ( // @[Xbar.scala 231:30]
    .clock(axi4xbar_clock),
    .reset(axi4xbar_reset),
    .auto_in_1_aw_ready(axi4xbar_auto_in_1_aw_ready),
    .auto_in_1_aw_valid(axi4xbar_auto_in_1_aw_valid),
    .auto_in_1_aw_bits_id(axi4xbar_auto_in_1_aw_bits_id),
    .auto_in_1_aw_bits_addr(axi4xbar_auto_in_1_aw_bits_addr),
    .auto_in_1_aw_bits_len(axi4xbar_auto_in_1_aw_bits_len),
    .auto_in_1_aw_bits_size(axi4xbar_auto_in_1_aw_bits_size),
    .auto_in_1_aw_bits_burst(axi4xbar_auto_in_1_aw_bits_burst),
    .auto_in_1_aw_bits_lock(axi4xbar_auto_in_1_aw_bits_lock),
    .auto_in_1_aw_bits_cache(axi4xbar_auto_in_1_aw_bits_cache),
    .auto_in_1_aw_bits_prot(axi4xbar_auto_in_1_aw_bits_prot),
    .auto_in_1_aw_bits_qos(axi4xbar_auto_in_1_aw_bits_qos),
    .auto_in_1_w_ready(axi4xbar_auto_in_1_w_ready),
    .auto_in_1_w_valid(axi4xbar_auto_in_1_w_valid),
    .auto_in_1_w_bits_data(axi4xbar_auto_in_1_w_bits_data),
    .auto_in_1_w_bits_strb(axi4xbar_auto_in_1_w_bits_strb),
    .auto_in_1_w_bits_last(axi4xbar_auto_in_1_w_bits_last),
    .auto_in_1_b_ready(axi4xbar_auto_in_1_b_ready),
    .auto_in_1_b_valid(axi4xbar_auto_in_1_b_valid),
    .auto_in_1_b_bits_id(axi4xbar_auto_in_1_b_bits_id),
    .auto_in_1_b_bits_resp(axi4xbar_auto_in_1_b_bits_resp),
    .auto_in_1_ar_ready(axi4xbar_auto_in_1_ar_ready),
    .auto_in_1_ar_valid(axi4xbar_auto_in_1_ar_valid),
    .auto_in_1_ar_bits_id(axi4xbar_auto_in_1_ar_bits_id),
    .auto_in_1_ar_bits_addr(axi4xbar_auto_in_1_ar_bits_addr),
    .auto_in_1_ar_bits_len(axi4xbar_auto_in_1_ar_bits_len),
    .auto_in_1_ar_bits_size(axi4xbar_auto_in_1_ar_bits_size),
    .auto_in_1_ar_bits_burst(axi4xbar_auto_in_1_ar_bits_burst),
    .auto_in_1_ar_bits_lock(axi4xbar_auto_in_1_ar_bits_lock),
    .auto_in_1_ar_bits_cache(axi4xbar_auto_in_1_ar_bits_cache),
    .auto_in_1_ar_bits_prot(axi4xbar_auto_in_1_ar_bits_prot),
    .auto_in_1_ar_bits_qos(axi4xbar_auto_in_1_ar_bits_qos),
    .auto_in_1_r_ready(axi4xbar_auto_in_1_r_ready),
    .auto_in_1_r_valid(axi4xbar_auto_in_1_r_valid),
    .auto_in_1_r_bits_id(axi4xbar_auto_in_1_r_bits_id),
    .auto_in_1_r_bits_data(axi4xbar_auto_in_1_r_bits_data),
    .auto_in_1_r_bits_resp(axi4xbar_auto_in_1_r_bits_resp),
    .auto_in_1_r_bits_last(axi4xbar_auto_in_1_r_bits_last),
    .auto_in_0_aw_ready(axi4xbar_auto_in_0_aw_ready),
    .auto_in_0_aw_valid(axi4xbar_auto_in_0_aw_valid),
    .auto_in_0_aw_bits_id(axi4xbar_auto_in_0_aw_bits_id),
    .auto_in_0_aw_bits_addr(axi4xbar_auto_in_0_aw_bits_addr),
    .auto_in_0_aw_bits_len(axi4xbar_auto_in_0_aw_bits_len),
    .auto_in_0_aw_bits_size(axi4xbar_auto_in_0_aw_bits_size),
    .auto_in_0_aw_bits_burst(axi4xbar_auto_in_0_aw_bits_burst),
    .auto_in_0_aw_bits_lock(axi4xbar_auto_in_0_aw_bits_lock),
    .auto_in_0_aw_bits_cache(axi4xbar_auto_in_0_aw_bits_cache),
    .auto_in_0_aw_bits_prot(axi4xbar_auto_in_0_aw_bits_prot),
    .auto_in_0_aw_bits_qos(axi4xbar_auto_in_0_aw_bits_qos),
    .auto_in_0_aw_bits_echo_tl_state_source(axi4xbar_auto_in_0_aw_bits_echo_tl_state_source),
    .auto_in_0_w_ready(axi4xbar_auto_in_0_w_ready),
    .auto_in_0_w_valid(axi4xbar_auto_in_0_w_valid),
    .auto_in_0_w_bits_data(axi4xbar_auto_in_0_w_bits_data),
    .auto_in_0_w_bits_strb(axi4xbar_auto_in_0_w_bits_strb),
    .auto_in_0_w_bits_last(axi4xbar_auto_in_0_w_bits_last),
    .auto_in_0_b_ready(axi4xbar_auto_in_0_b_ready),
    .auto_in_0_b_valid(axi4xbar_auto_in_0_b_valid),
    .auto_in_0_b_bits_id(axi4xbar_auto_in_0_b_bits_id),
    .auto_in_0_b_bits_echo_tl_state_source(axi4xbar_auto_in_0_b_bits_echo_tl_state_source),
    .auto_in_0_ar_ready(axi4xbar_auto_in_0_ar_ready),
    .auto_in_0_ar_valid(axi4xbar_auto_in_0_ar_valid),
    .auto_in_0_ar_bits_id(axi4xbar_auto_in_0_ar_bits_id),
    .auto_in_0_ar_bits_addr(axi4xbar_auto_in_0_ar_bits_addr),
    .auto_in_0_ar_bits_len(axi4xbar_auto_in_0_ar_bits_len),
    .auto_in_0_ar_bits_size(axi4xbar_auto_in_0_ar_bits_size),
    .auto_in_0_ar_bits_burst(axi4xbar_auto_in_0_ar_bits_burst),
    .auto_in_0_ar_bits_lock(axi4xbar_auto_in_0_ar_bits_lock),
    .auto_in_0_ar_bits_cache(axi4xbar_auto_in_0_ar_bits_cache),
    .auto_in_0_ar_bits_prot(axi4xbar_auto_in_0_ar_bits_prot),
    .auto_in_0_ar_bits_qos(axi4xbar_auto_in_0_ar_bits_qos),
    .auto_in_0_ar_bits_echo_tl_state_source(axi4xbar_auto_in_0_ar_bits_echo_tl_state_source),
    .auto_in_0_r_ready(axi4xbar_auto_in_0_r_ready),
    .auto_in_0_r_valid(axi4xbar_auto_in_0_r_valid),
    .auto_in_0_r_bits_id(axi4xbar_auto_in_0_r_bits_id),
    .auto_in_0_r_bits_data(axi4xbar_auto_in_0_r_bits_data),
    .auto_in_0_r_bits_echo_tl_state_source(axi4xbar_auto_in_0_r_bits_echo_tl_state_source),
    .auto_in_0_r_bits_last(axi4xbar_auto_in_0_r_bits_last),
    .auto_out_aw_ready(axi4xbar_auto_out_aw_ready),
    .auto_out_aw_valid(axi4xbar_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4xbar_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4xbar_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4xbar_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4xbar_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(axi4xbar_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(axi4xbar_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(axi4xbar_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(axi4xbar_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(axi4xbar_auto_out_aw_bits_qos),
    .auto_out_aw_bits_echo_tl_state_source(axi4xbar_auto_out_aw_bits_echo_tl_state_source),
    .auto_out_w_ready(axi4xbar_auto_out_w_ready),
    .auto_out_w_valid(axi4xbar_auto_out_w_valid),
    .auto_out_w_bits_data(axi4xbar_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4xbar_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4xbar_auto_out_w_bits_last),
    .auto_out_b_ready(axi4xbar_auto_out_b_ready),
    .auto_out_b_valid(axi4xbar_auto_out_b_valid),
    .auto_out_b_bits_id(axi4xbar_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4xbar_auto_out_b_bits_resp),
    .auto_out_b_bits_echo_tl_state_source(axi4xbar_auto_out_b_bits_echo_tl_state_source),
    .auto_out_ar_ready(axi4xbar_auto_out_ar_ready),
    .auto_out_ar_valid(axi4xbar_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4xbar_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4xbar_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4xbar_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4xbar_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(axi4xbar_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(axi4xbar_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(axi4xbar_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(axi4xbar_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(axi4xbar_auto_out_ar_bits_qos),
    .auto_out_ar_bits_echo_tl_state_source(axi4xbar_auto_out_ar_bits_echo_tl_state_source),
    .auto_out_r_ready(axi4xbar_auto_out_r_ready),
    .auto_out_r_valid(axi4xbar_auto_out_r_valid),
    .auto_out_r_bits_id(axi4xbar_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4xbar_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4xbar_auto_out_r_bits_resp),
    .auto_out_r_bits_echo_tl_state_source(axi4xbar_auto_out_r_bits_echo_tl_state_source),
    .auto_out_r_bits_last(axi4xbar_auto_out_r_bits_last)
  );
  AXI4Xbar_1 axi4xbar_1 ( // @[Xbar.scala 231:30]
    .clock(axi4xbar_1_clock),
    .reset(axi4xbar_1_reset),
    .auto_in_aw_ready(axi4xbar_1_auto_in_aw_ready),
    .auto_in_aw_valid(axi4xbar_1_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4xbar_1_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4xbar_1_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4xbar_1_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4xbar_1_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axi4xbar_1_auto_in_aw_bits_burst),
    .auto_in_aw_bits_lock(axi4xbar_1_auto_in_aw_bits_lock),
    .auto_in_aw_bits_cache(axi4xbar_1_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(axi4xbar_1_auto_in_aw_bits_prot),
    .auto_in_aw_bits_qos(axi4xbar_1_auto_in_aw_bits_qos),
    .auto_in_w_ready(axi4xbar_1_auto_in_w_ready),
    .auto_in_w_valid(axi4xbar_1_auto_in_w_valid),
    .auto_in_w_bits_data(axi4xbar_1_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4xbar_1_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4xbar_1_auto_in_w_bits_last),
    .auto_in_b_ready(axi4xbar_1_auto_in_b_ready),
    .auto_in_b_valid(axi4xbar_1_auto_in_b_valid),
    .auto_in_b_bits_id(axi4xbar_1_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4xbar_1_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4xbar_1_auto_in_ar_ready),
    .auto_in_ar_valid(axi4xbar_1_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4xbar_1_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4xbar_1_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4xbar_1_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4xbar_1_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axi4xbar_1_auto_in_ar_bits_burst),
    .auto_in_ar_bits_lock(axi4xbar_1_auto_in_ar_bits_lock),
    .auto_in_ar_bits_cache(axi4xbar_1_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(axi4xbar_1_auto_in_ar_bits_prot),
    .auto_in_ar_bits_qos(axi4xbar_1_auto_in_ar_bits_qos),
    .auto_in_r_ready(axi4xbar_1_auto_in_r_ready),
    .auto_in_r_valid(axi4xbar_1_auto_in_r_valid),
    .auto_in_r_bits_id(axi4xbar_1_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4xbar_1_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4xbar_1_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4xbar_1_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4xbar_1_auto_out_aw_ready),
    .auto_out_aw_valid(axi4xbar_1_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4xbar_1_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4xbar_1_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4xbar_1_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4xbar_1_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(axi4xbar_1_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(axi4xbar_1_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(axi4xbar_1_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(axi4xbar_1_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(axi4xbar_1_auto_out_aw_bits_qos),
    .auto_out_w_ready(axi4xbar_1_auto_out_w_ready),
    .auto_out_w_valid(axi4xbar_1_auto_out_w_valid),
    .auto_out_w_bits_data(axi4xbar_1_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4xbar_1_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4xbar_1_auto_out_w_bits_last),
    .auto_out_b_ready(axi4xbar_1_auto_out_b_ready),
    .auto_out_b_valid(axi4xbar_1_auto_out_b_valid),
    .auto_out_b_bits_id(axi4xbar_1_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4xbar_1_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4xbar_1_auto_out_ar_ready),
    .auto_out_ar_valid(axi4xbar_1_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4xbar_1_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4xbar_1_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4xbar_1_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4xbar_1_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(axi4xbar_1_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(axi4xbar_1_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(axi4xbar_1_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(axi4xbar_1_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(axi4xbar_1_auto_out_ar_bits_qos),
    .auto_out_r_ready(axi4xbar_1_auto_out_r_ready),
    .auto_out_r_valid(axi4xbar_1_auto_out_r_valid),
    .auto_out_r_bits_id(axi4xbar_1_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4xbar_1_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4xbar_1_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4xbar_1_auto_out_r_bits_last)
  );
  AXI4Buffer_2 axi4buf_2 ( // @[Buffer.scala 63:29]
    .clock(axi4buf_2_clock),
    .reset(axi4buf_2_reset),
    .auto_in_aw_ready(axi4buf_2_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_2_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_2_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_2_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4buf_2_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4buf_2_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axi4buf_2_auto_in_aw_bits_burst),
    .auto_in_aw_bits_lock(axi4buf_2_auto_in_aw_bits_lock),
    .auto_in_aw_bits_cache(axi4buf_2_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(axi4buf_2_auto_in_aw_bits_prot),
    .auto_in_aw_bits_qos(axi4buf_2_auto_in_aw_bits_qos),
    .auto_in_w_ready(axi4buf_2_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_2_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_2_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_2_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_2_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_2_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_2_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_2_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_2_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_2_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_2_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_2_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_2_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4buf_2_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4buf_2_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axi4buf_2_auto_in_ar_bits_burst),
    .auto_in_ar_bits_lock(axi4buf_2_auto_in_ar_bits_lock),
    .auto_in_ar_bits_cache(axi4buf_2_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(axi4buf_2_auto_in_ar_bits_prot),
    .auto_in_ar_bits_qos(axi4buf_2_auto_in_ar_bits_qos),
    .auto_in_r_ready(axi4buf_2_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_2_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_2_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_2_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_2_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_2_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_2_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_2_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_2_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_2_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4buf_2_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4buf_2_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(axi4buf_2_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(axi4buf_2_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(axi4buf_2_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(axi4buf_2_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(axi4buf_2_auto_out_aw_bits_qos),
    .auto_out_w_ready(axi4buf_2_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_2_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_2_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_2_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_2_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_2_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_2_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_2_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_2_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_2_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_2_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_2_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_2_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4buf_2_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4buf_2_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(axi4buf_2_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(axi4buf_2_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(axi4buf_2_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(axi4buf_2_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(axi4buf_2_auto_out_ar_bits_qos),
    .auto_out_r_ready(axi4buf_2_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_2_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_2_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_2_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_2_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_2_auto_out_r_bits_last)
  );
  AXI4Buffer_2 axi4buf_3 ( // @[Buffer.scala 63:29]
    .clock(axi4buf_3_clock),
    .reset(axi4buf_3_reset),
    .auto_in_aw_ready(axi4buf_3_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_3_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_3_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_3_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4buf_3_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4buf_3_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axi4buf_3_auto_in_aw_bits_burst),
    .auto_in_aw_bits_lock(axi4buf_3_auto_in_aw_bits_lock),
    .auto_in_aw_bits_cache(axi4buf_3_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(axi4buf_3_auto_in_aw_bits_prot),
    .auto_in_aw_bits_qos(axi4buf_3_auto_in_aw_bits_qos),
    .auto_in_w_ready(axi4buf_3_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_3_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_3_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_3_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_3_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_3_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_3_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_3_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_3_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_3_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_3_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_3_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_3_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4buf_3_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4buf_3_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axi4buf_3_auto_in_ar_bits_burst),
    .auto_in_ar_bits_lock(axi4buf_3_auto_in_ar_bits_lock),
    .auto_in_ar_bits_cache(axi4buf_3_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(axi4buf_3_auto_in_ar_bits_prot),
    .auto_in_ar_bits_qos(axi4buf_3_auto_in_ar_bits_qos),
    .auto_in_r_ready(axi4buf_3_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_3_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_3_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_3_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_3_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_3_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_3_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_3_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_3_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_3_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4buf_3_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4buf_3_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(axi4buf_3_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(axi4buf_3_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(axi4buf_3_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(axi4buf_3_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(axi4buf_3_auto_out_aw_bits_qos),
    .auto_out_w_ready(axi4buf_3_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_3_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_3_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_3_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_3_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_3_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_3_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_3_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_3_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_3_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_3_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_3_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_3_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4buf_3_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4buf_3_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(axi4buf_3_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(axi4buf_3_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(axi4buf_3_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(axi4buf_3_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(axi4buf_3_auto_out_ar_bits_qos),
    .auto_out_r_ready(axi4buf_3_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_3_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_3_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_3_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_3_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_3_auto_out_r_bits_last)
  );
  AXI4UserYanker axi4yank ( // @[UserYanker.scala 108:30]
    .clock(axi4yank_clock),
    .reset(axi4yank_reset),
    .auto_in_aw_ready(axi4yank_auto_in_aw_ready),
    .auto_in_aw_valid(axi4yank_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4yank_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4yank_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4yank_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4yank_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axi4yank_auto_in_aw_bits_burst),
    .auto_in_aw_bits_lock(axi4yank_auto_in_aw_bits_lock),
    .auto_in_aw_bits_cache(axi4yank_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(axi4yank_auto_in_aw_bits_prot),
    .auto_in_aw_bits_qos(axi4yank_auto_in_aw_bits_qos),
    .auto_in_aw_bits_echo_tl_state_source(axi4yank_auto_in_aw_bits_echo_tl_state_source),
    .auto_in_aw_bits_echo_extra_id(axi4yank_auto_in_aw_bits_echo_extra_id),
    .auto_in_w_ready(axi4yank_auto_in_w_ready),
    .auto_in_w_valid(axi4yank_auto_in_w_valid),
    .auto_in_w_bits_data(axi4yank_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4yank_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4yank_auto_in_w_bits_last),
    .auto_in_b_ready(axi4yank_auto_in_b_ready),
    .auto_in_b_valid(axi4yank_auto_in_b_valid),
    .auto_in_b_bits_id(axi4yank_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4yank_auto_in_b_bits_resp),
    .auto_in_b_bits_echo_tl_state_source(axi4yank_auto_in_b_bits_echo_tl_state_source),
    .auto_in_b_bits_echo_extra_id(axi4yank_auto_in_b_bits_echo_extra_id),
    .auto_in_ar_ready(axi4yank_auto_in_ar_ready),
    .auto_in_ar_valid(axi4yank_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4yank_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4yank_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4yank_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4yank_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axi4yank_auto_in_ar_bits_burst),
    .auto_in_ar_bits_lock(axi4yank_auto_in_ar_bits_lock),
    .auto_in_ar_bits_cache(axi4yank_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(axi4yank_auto_in_ar_bits_prot),
    .auto_in_ar_bits_qos(axi4yank_auto_in_ar_bits_qos),
    .auto_in_ar_bits_echo_tl_state_source(axi4yank_auto_in_ar_bits_echo_tl_state_source),
    .auto_in_ar_bits_echo_extra_id(axi4yank_auto_in_ar_bits_echo_extra_id),
    .auto_in_r_ready(axi4yank_auto_in_r_ready),
    .auto_in_r_valid(axi4yank_auto_in_r_valid),
    .auto_in_r_bits_id(axi4yank_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4yank_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4yank_auto_in_r_bits_resp),
    .auto_in_r_bits_echo_tl_state_source(axi4yank_auto_in_r_bits_echo_tl_state_source),
    .auto_in_r_bits_echo_extra_id(axi4yank_auto_in_r_bits_echo_extra_id),
    .auto_in_r_bits_last(axi4yank_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4yank_auto_out_aw_ready),
    .auto_out_aw_valid(axi4yank_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4yank_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4yank_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4yank_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4yank_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(axi4yank_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(axi4yank_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(axi4yank_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(axi4yank_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(axi4yank_auto_out_aw_bits_qos),
    .auto_out_w_ready(axi4yank_auto_out_w_ready),
    .auto_out_w_valid(axi4yank_auto_out_w_valid),
    .auto_out_w_bits_data(axi4yank_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4yank_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4yank_auto_out_w_bits_last),
    .auto_out_b_ready(axi4yank_auto_out_b_ready),
    .auto_out_b_valid(axi4yank_auto_out_b_valid),
    .auto_out_b_bits_id(axi4yank_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4yank_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4yank_auto_out_ar_ready),
    .auto_out_ar_valid(axi4yank_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4yank_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4yank_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4yank_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4yank_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(axi4yank_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(axi4yank_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(axi4yank_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(axi4yank_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(axi4yank_auto_out_ar_bits_qos),
    .auto_out_r_ready(axi4yank_auto_out_r_ready),
    .auto_out_r_valid(axi4yank_auto_out_r_valid),
    .auto_out_r_bits_id(axi4yank_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4yank_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4yank_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4yank_auto_out_r_bits_last)
  );
  AXI4Buffer_4 axi4buf_4 ( // @[Buffer.scala 63:29]
    .clock(axi4buf_4_clock),
    .reset(axi4buf_4_reset),
    .auto_in_aw_ready(axi4buf_4_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_4_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_4_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_4_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4buf_4_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4buf_4_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axi4buf_4_auto_in_aw_bits_burst),
    .auto_in_aw_bits_lock(axi4buf_4_auto_in_aw_bits_lock),
    .auto_in_aw_bits_cache(axi4buf_4_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(axi4buf_4_auto_in_aw_bits_prot),
    .auto_in_aw_bits_qos(axi4buf_4_auto_in_aw_bits_qos),
    .auto_in_aw_bits_echo_tl_state_source(axi4buf_4_auto_in_aw_bits_echo_tl_state_source),
    .auto_in_aw_bits_echo_extra_id(axi4buf_4_auto_in_aw_bits_echo_extra_id),
    .auto_in_w_ready(axi4buf_4_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_4_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_4_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_4_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_4_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_4_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_4_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_4_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_4_auto_in_b_bits_resp),
    .auto_in_b_bits_echo_tl_state_source(axi4buf_4_auto_in_b_bits_echo_tl_state_source),
    .auto_in_b_bits_echo_extra_id(axi4buf_4_auto_in_b_bits_echo_extra_id),
    .auto_in_ar_ready(axi4buf_4_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_4_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_4_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_4_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4buf_4_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4buf_4_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axi4buf_4_auto_in_ar_bits_burst),
    .auto_in_ar_bits_lock(axi4buf_4_auto_in_ar_bits_lock),
    .auto_in_ar_bits_cache(axi4buf_4_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(axi4buf_4_auto_in_ar_bits_prot),
    .auto_in_ar_bits_qos(axi4buf_4_auto_in_ar_bits_qos),
    .auto_in_ar_bits_echo_tl_state_source(axi4buf_4_auto_in_ar_bits_echo_tl_state_source),
    .auto_in_ar_bits_echo_extra_id(axi4buf_4_auto_in_ar_bits_echo_extra_id),
    .auto_in_r_ready(axi4buf_4_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_4_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_4_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_4_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_4_auto_in_r_bits_resp),
    .auto_in_r_bits_echo_tl_state_source(axi4buf_4_auto_in_r_bits_echo_tl_state_source),
    .auto_in_r_bits_echo_extra_id(axi4buf_4_auto_in_r_bits_echo_extra_id),
    .auto_in_r_bits_last(axi4buf_4_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_4_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_4_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_4_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_4_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4buf_4_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4buf_4_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(axi4buf_4_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(axi4buf_4_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(axi4buf_4_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(axi4buf_4_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(axi4buf_4_auto_out_aw_bits_qos),
    .auto_out_aw_bits_echo_tl_state_source(axi4buf_4_auto_out_aw_bits_echo_tl_state_source),
    .auto_out_aw_bits_echo_extra_id(axi4buf_4_auto_out_aw_bits_echo_extra_id),
    .auto_out_w_ready(axi4buf_4_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_4_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_4_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_4_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_4_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_4_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_4_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_4_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_4_auto_out_b_bits_resp),
    .auto_out_b_bits_echo_tl_state_source(axi4buf_4_auto_out_b_bits_echo_tl_state_source),
    .auto_out_b_bits_echo_extra_id(axi4buf_4_auto_out_b_bits_echo_extra_id),
    .auto_out_ar_ready(axi4buf_4_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_4_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_4_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_4_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4buf_4_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4buf_4_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(axi4buf_4_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(axi4buf_4_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(axi4buf_4_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(axi4buf_4_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(axi4buf_4_auto_out_ar_bits_qos),
    .auto_out_ar_bits_echo_tl_state_source(axi4buf_4_auto_out_ar_bits_echo_tl_state_source),
    .auto_out_ar_bits_echo_extra_id(axi4buf_4_auto_out_ar_bits_echo_extra_id),
    .auto_out_r_ready(axi4buf_4_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_4_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_4_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_4_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_4_auto_out_r_bits_resp),
    .auto_out_r_bits_echo_tl_state_source(axi4buf_4_auto_out_r_bits_echo_tl_state_source),
    .auto_out_r_bits_echo_extra_id(axi4buf_4_auto_out_r_bits_echo_extra_id),
    .auto_out_r_bits_last(axi4buf_4_auto_out_r_bits_last)
  );
  AXI4IdIndexer axi4index ( // @[IdIndexer.scala 94:31]
    .auto_in_aw_ready(axi4index_auto_in_aw_ready),
    .auto_in_aw_valid(axi4index_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4index_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4index_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4index_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4index_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axi4index_auto_in_aw_bits_burst),
    .auto_in_aw_bits_lock(axi4index_auto_in_aw_bits_lock),
    .auto_in_aw_bits_cache(axi4index_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(axi4index_auto_in_aw_bits_prot),
    .auto_in_aw_bits_qos(axi4index_auto_in_aw_bits_qos),
    .auto_in_aw_bits_echo_tl_state_source(axi4index_auto_in_aw_bits_echo_tl_state_source),
    .auto_in_w_ready(axi4index_auto_in_w_ready),
    .auto_in_w_valid(axi4index_auto_in_w_valid),
    .auto_in_w_bits_data(axi4index_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4index_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4index_auto_in_w_bits_last),
    .auto_in_b_ready(axi4index_auto_in_b_ready),
    .auto_in_b_valid(axi4index_auto_in_b_valid),
    .auto_in_b_bits_id(axi4index_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4index_auto_in_b_bits_resp),
    .auto_in_b_bits_echo_tl_state_source(axi4index_auto_in_b_bits_echo_tl_state_source),
    .auto_in_ar_ready(axi4index_auto_in_ar_ready),
    .auto_in_ar_valid(axi4index_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4index_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4index_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4index_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4index_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axi4index_auto_in_ar_bits_burst),
    .auto_in_ar_bits_lock(axi4index_auto_in_ar_bits_lock),
    .auto_in_ar_bits_cache(axi4index_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(axi4index_auto_in_ar_bits_prot),
    .auto_in_ar_bits_qos(axi4index_auto_in_ar_bits_qos),
    .auto_in_ar_bits_echo_tl_state_source(axi4index_auto_in_ar_bits_echo_tl_state_source),
    .auto_in_r_ready(axi4index_auto_in_r_ready),
    .auto_in_r_valid(axi4index_auto_in_r_valid),
    .auto_in_r_bits_id(axi4index_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4index_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4index_auto_in_r_bits_resp),
    .auto_in_r_bits_echo_tl_state_source(axi4index_auto_in_r_bits_echo_tl_state_source),
    .auto_in_r_bits_last(axi4index_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4index_auto_out_aw_ready),
    .auto_out_aw_valid(axi4index_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4index_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4index_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4index_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4index_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(axi4index_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(axi4index_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(axi4index_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(axi4index_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(axi4index_auto_out_aw_bits_qos),
    .auto_out_aw_bits_echo_tl_state_source(axi4index_auto_out_aw_bits_echo_tl_state_source),
    .auto_out_aw_bits_echo_extra_id(axi4index_auto_out_aw_bits_echo_extra_id),
    .auto_out_w_ready(axi4index_auto_out_w_ready),
    .auto_out_w_valid(axi4index_auto_out_w_valid),
    .auto_out_w_bits_data(axi4index_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4index_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4index_auto_out_w_bits_last),
    .auto_out_b_ready(axi4index_auto_out_b_ready),
    .auto_out_b_valid(axi4index_auto_out_b_valid),
    .auto_out_b_bits_id(axi4index_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4index_auto_out_b_bits_resp),
    .auto_out_b_bits_echo_tl_state_source(axi4index_auto_out_b_bits_echo_tl_state_source),
    .auto_out_b_bits_echo_extra_id(axi4index_auto_out_b_bits_echo_extra_id),
    .auto_out_ar_ready(axi4index_auto_out_ar_ready),
    .auto_out_ar_valid(axi4index_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4index_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4index_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4index_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4index_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(axi4index_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(axi4index_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(axi4index_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(axi4index_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(axi4index_auto_out_ar_bits_qos),
    .auto_out_ar_bits_echo_tl_state_source(axi4index_auto_out_ar_bits_echo_tl_state_source),
    .auto_out_ar_bits_echo_extra_id(axi4index_auto_out_ar_bits_echo_extra_id),
    .auto_out_r_ready(axi4index_auto_out_r_ready),
    .auto_out_r_valid(axi4index_auto_out_r_valid),
    .auto_out_r_bits_id(axi4index_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4index_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4index_auto_out_r_bits_resp),
    .auto_out_r_bits_echo_tl_state_source(axi4index_auto_out_r_bits_echo_tl_state_source),
    .auto_out_r_bits_echo_extra_id(axi4index_auto_out_r_bits_echo_extra_id),
    .auto_out_r_bits_last(axi4index_auto_out_r_bits_last)
  );
  AXI4Buffer_5 axi4buf_5 ( // @[Buffer.scala 63:29]
    .clock(axi4buf_5_clock),
    .reset(axi4buf_5_reset),
    .auto_in_aw_ready(axi4buf_5_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_5_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_5_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_5_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4buf_5_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4buf_5_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axi4buf_5_auto_in_aw_bits_burst),
    .auto_in_aw_bits_lock(axi4buf_5_auto_in_aw_bits_lock),
    .auto_in_aw_bits_cache(axi4buf_5_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(axi4buf_5_auto_in_aw_bits_prot),
    .auto_in_aw_bits_qos(axi4buf_5_auto_in_aw_bits_qos),
    .auto_in_aw_bits_echo_tl_state_source(axi4buf_5_auto_in_aw_bits_echo_tl_state_source),
    .auto_in_w_ready(axi4buf_5_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_5_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_5_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_5_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_5_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_5_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_5_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_5_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_5_auto_in_b_bits_resp),
    .auto_in_b_bits_echo_tl_state_source(axi4buf_5_auto_in_b_bits_echo_tl_state_source),
    .auto_in_ar_ready(axi4buf_5_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_5_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_5_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_5_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4buf_5_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4buf_5_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axi4buf_5_auto_in_ar_bits_burst),
    .auto_in_ar_bits_lock(axi4buf_5_auto_in_ar_bits_lock),
    .auto_in_ar_bits_cache(axi4buf_5_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(axi4buf_5_auto_in_ar_bits_prot),
    .auto_in_ar_bits_qos(axi4buf_5_auto_in_ar_bits_qos),
    .auto_in_ar_bits_echo_tl_state_source(axi4buf_5_auto_in_ar_bits_echo_tl_state_source),
    .auto_in_r_ready(axi4buf_5_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_5_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_5_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_5_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_5_auto_in_r_bits_resp),
    .auto_in_r_bits_echo_tl_state_source(axi4buf_5_auto_in_r_bits_echo_tl_state_source),
    .auto_in_r_bits_last(axi4buf_5_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_5_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_5_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_5_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_5_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4buf_5_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4buf_5_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(axi4buf_5_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(axi4buf_5_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(axi4buf_5_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(axi4buf_5_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(axi4buf_5_auto_out_aw_bits_qos),
    .auto_out_aw_bits_echo_tl_state_source(axi4buf_5_auto_out_aw_bits_echo_tl_state_source),
    .auto_out_w_ready(axi4buf_5_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_5_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_5_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_5_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_5_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_5_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_5_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_5_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_5_auto_out_b_bits_resp),
    .auto_out_b_bits_echo_tl_state_source(axi4buf_5_auto_out_b_bits_echo_tl_state_source),
    .auto_out_ar_ready(axi4buf_5_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_5_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_5_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_5_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4buf_5_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4buf_5_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(axi4buf_5_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(axi4buf_5_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(axi4buf_5_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(axi4buf_5_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(axi4buf_5_auto_out_ar_bits_qos),
    .auto_out_ar_bits_echo_tl_state_source(axi4buf_5_auto_out_ar_bits_echo_tl_state_source),
    .auto_out_r_ready(axi4buf_5_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_5_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_5_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_5_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_5_auto_out_r_bits_resp),
    .auto_out_r_bits_echo_tl_state_source(axi4buf_5_auto_out_r_bits_echo_tl_state_source),
    .auto_out_r_bits_last(axi4buf_5_auto_out_r_bits_last)
  );
  AXILHub cmd_resp_axilhub ( // @[ComposerTop.scala 134:36]
    .clock(cmd_resp_axilhub_clock),
    .reset(cmd_resp_axilhub_reset),
    .auto_in_aw_ready(cmd_resp_axilhub_auto_in_aw_ready),
    .auto_in_aw_valid(cmd_resp_axilhub_auto_in_aw_valid),
    .auto_in_aw_bits_id(cmd_resp_axilhub_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(cmd_resp_axilhub_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(cmd_resp_axilhub_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(cmd_resp_axilhub_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(cmd_resp_axilhub_auto_in_aw_bits_burst),
    .auto_in_w_ready(cmd_resp_axilhub_auto_in_w_ready),
    .auto_in_w_valid(cmd_resp_axilhub_auto_in_w_valid),
    .auto_in_w_bits_data(cmd_resp_axilhub_auto_in_w_bits_data),
    .auto_in_w_bits_last(cmd_resp_axilhub_auto_in_w_bits_last),
    .auto_in_b_ready(cmd_resp_axilhub_auto_in_b_ready),
    .auto_in_b_valid(cmd_resp_axilhub_auto_in_b_valid),
    .auto_in_b_bits_id(cmd_resp_axilhub_auto_in_b_bits_id),
    .auto_in_b_bits_resp(cmd_resp_axilhub_auto_in_b_bits_resp),
    .auto_in_ar_ready(cmd_resp_axilhub_auto_in_ar_ready),
    .auto_in_ar_valid(cmd_resp_axilhub_auto_in_ar_valid),
    .auto_in_ar_bits_id(cmd_resp_axilhub_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(cmd_resp_axilhub_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(cmd_resp_axilhub_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(cmd_resp_axilhub_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(cmd_resp_axilhub_auto_in_ar_bits_burst),
    .auto_in_r_ready(cmd_resp_axilhub_auto_in_r_ready),
    .auto_in_r_valid(cmd_resp_axilhub_auto_in_r_valid),
    .auto_in_r_bits_id(cmd_resp_axilhub_auto_in_r_bits_id),
    .auto_in_r_bits_data(cmd_resp_axilhub_auto_in_r_bits_data),
    .auto_in_r_bits_resp(cmd_resp_axilhub_auto_in_r_bits_resp),
    .auto_in_r_bits_last(cmd_resp_axilhub_auto_in_r_bits_last),
    .io_rocc_in_ready(cmd_resp_axilhub_io_rocc_in_ready),
    .io_rocc_in_valid(cmd_resp_axilhub_io_rocc_in_valid),
    .io_rocc_in_bits_inst_funct(cmd_resp_axilhub_io_rocc_in_bits_inst_funct),
    .io_rocc_in_bits_inst_rs2(cmd_resp_axilhub_io_rocc_in_bits_inst_rs2),
    .io_rocc_in_bits_inst_rs1(cmd_resp_axilhub_io_rocc_in_bits_inst_rs1),
    .io_rocc_in_bits_inst_opcode(cmd_resp_axilhub_io_rocc_in_bits_inst_opcode),
    .io_rocc_in_bits_rs1(cmd_resp_axilhub_io_rocc_in_bits_rs1),
    .io_rocc_in_bits_rs2(cmd_resp_axilhub_io_rocc_in_bits_rs2),
    .io_rocc_out_ready(cmd_resp_axilhub_io_rocc_out_ready),
    .io_rocc_out_valid(cmd_resp_axilhub_io_rocc_out_valid),
    .io_rocc_out_bits_rd(cmd_resp_axilhub_io_rocc_out_bits_rd),
    .io_rocc_out_bits_data(cmd_resp_axilhub_io_rocc_out_bits_data)
  );
  AXI4Buffer_6 axi4buf_6 ( // @[Buffer.scala 63:29]
    .clock(axi4buf_6_clock),
    .reset(axi4buf_6_reset),
    .auto_in_aw_ready(axi4buf_6_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_6_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_6_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_6_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4buf_6_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4buf_6_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axi4buf_6_auto_in_aw_bits_burst),
    .auto_in_w_ready(axi4buf_6_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_6_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_6_auto_in_w_bits_data),
    .auto_in_w_bits_last(axi4buf_6_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_6_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_6_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_6_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_6_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_6_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_6_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_6_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_6_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4buf_6_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4buf_6_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axi4buf_6_auto_in_ar_bits_burst),
    .auto_in_r_ready(axi4buf_6_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_6_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_6_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_6_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_6_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_6_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_6_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_6_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_6_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_6_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4buf_6_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4buf_6_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(axi4buf_6_auto_out_aw_bits_burst),
    .auto_out_w_ready(axi4buf_6_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_6_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_6_auto_out_w_bits_data),
    .auto_out_w_bits_last(axi4buf_6_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_6_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_6_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_6_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_6_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_6_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_6_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_6_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_6_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4buf_6_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4buf_6_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(axi4buf_6_auto_out_ar_bits_burst),
    .auto_out_r_ready(axi4buf_6_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_6_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_6_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_6_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_6_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_6_auto_out_r_bits_last)
  );
  assign S00_AXI_awready = axi4buf_6_auto_in_aw_ready; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign S00_AXI_wready = axi4buf_6_auto_in_w_ready; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign S00_AXI_bid = axi4buf_6_auto_in_b_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign S00_AXI_bresp = axi4buf_6_auto_in_b_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign S00_AXI_bvalid = axi4buf_6_auto_in_b_valid; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign S00_AXI_arready = axi4buf_6_auto_in_ar_ready; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign S00_AXI_rid = axi4buf_6_auto_in_r_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign S00_AXI_rdata = axi4buf_6_auto_in_r_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign S00_AXI_rresp = axi4buf_6_auto_in_r_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign S00_AXI_rlast = axi4buf_6_auto_in_r_bits_last; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign S00_AXI_rvalid = axi4buf_6_auto_in_r_valid; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign M00_AXI_awid = axi4buf_3_auto_out_aw_bits_id; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_awaddr = axi4buf_3_auto_out_aw_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_awlen = axi4buf_3_auto_out_aw_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_awsize = axi4buf_3_auto_out_aw_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_awburst = axi4buf_3_auto_out_aw_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_awlock = axi4buf_3_auto_out_aw_bits_lock; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_awcache = axi4buf_3_auto_out_aw_bits_cache; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_awprot = axi4buf_3_auto_out_aw_bits_prot; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_awregion = 4'h0; // @[AXI4Compat.scala 90:21]
  assign M00_AXI_awqos = axi4buf_3_auto_out_aw_bits_qos; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_awvalid = axi4buf_3_auto_out_aw_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_wdata = axi4buf_3_auto_out_w_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_wstrb = axi4buf_3_auto_out_w_bits_strb; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_wlast = axi4buf_3_auto_out_w_bits_last; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_wvalid = axi4buf_3_auto_out_w_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_bready = axi4buf_3_auto_out_b_ready; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_arid = axi4buf_3_auto_out_ar_bits_id; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_araddr = axi4buf_3_auto_out_ar_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_arlen = axi4buf_3_auto_out_ar_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_arsize = axi4buf_3_auto_out_ar_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_arburst = axi4buf_3_auto_out_ar_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_arlock = axi4buf_3_auto_out_ar_bits_lock; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_arcache = axi4buf_3_auto_out_ar_bits_cache; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_arprot = axi4buf_3_auto_out_ar_bits_prot; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_arregion = 4'h0; // @[AXI4Compat.scala 71:21]
  assign M00_AXI_arqos = axi4buf_3_auto_out_ar_bits_qos; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_arvalid = axi4buf_3_auto_out_ar_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign M00_AXI_rready = axi4buf_3_auto_out_r_ready; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign dma_awready = axi4buf_2_auto_in_aw_ready; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign dma_wready = axi4buf_2_auto_in_w_ready; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign dma_bid = axi4buf_2_auto_in_b_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign dma_bresp = axi4buf_2_auto_in_b_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign dma_bvalid = axi4buf_2_auto_in_b_valid; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign dma_arready = axi4buf_2_auto_in_ar_ready; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign dma_rid = axi4buf_2_auto_in_r_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign dma_rdata = axi4buf_2_auto_in_r_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign dma_rresp = axi4buf_2_auto_in_r_bits_resp; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign dma_rlast = axi4buf_2_auto_in_r_bits_last; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign dma_rvalid = axi4buf_2_auto_in_r_valid; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign acc_clock = clock;
  assign acc_reset = reset;
  assign acc_auto_mem_out_a_ready = tl2axi4_auto_in_a_ready; // @[LazyModule.scala 355:16]
  assign acc_auto_mem_out_d_valid = tl2axi4_auto_in_d_valid; // @[LazyModule.scala 355:16]
  assign acc_auto_mem_out_d_bits_source = tl2axi4_auto_in_d_bits_source; // @[LazyModule.scala 355:16]
  assign acc_auto_mem_out_d_bits_data = tl2axi4_auto_in_d_bits_data; // @[LazyModule.scala 355:16]
  assign acc_io_cmd_valid = cmd_resp_axilhub_io_rocc_in_valid; // @[ComposerTop.scala 148:21]
  assign acc_io_cmd_bits_inst_funct = cmd_resp_axilhub_io_rocc_in_bits_inst_funct; // @[ComposerTop.scala 148:21]
  assign acc_io_cmd_bits_inst_rs2 = cmd_resp_axilhub_io_rocc_in_bits_inst_rs2; // @[ComposerTop.scala 148:21]
  assign acc_io_cmd_bits_inst_rs1 = cmd_resp_axilhub_io_rocc_in_bits_inst_rs1; // @[ComposerTop.scala 148:21]
  assign acc_io_cmd_bits_inst_opcode = cmd_resp_axilhub_io_rocc_in_bits_inst_opcode; // @[ComposerTop.scala 148:21]
  assign acc_io_cmd_bits_rs1 = cmd_resp_axilhub_io_rocc_in_bits_rs1; // @[ComposerTop.scala 148:21]
  assign acc_io_cmd_bits_rs2 = cmd_resp_axilhub_io_rocc_in_bits_rs2; // @[ComposerTop.scala 148:21]
  assign acc_io_resp_ready = cmd_resp_axilhub_io_rocc_out_ready; // @[ComposerTop.scala 149:31]
  assign axi4buf_clock = clock;
  assign axi4buf_reset = reset;
  assign axi4buf_auto_in_aw_valid = axi4buf_1_auto_out_aw_valid; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_aw_bits_id = axi4buf_1_auto_out_aw_bits_id; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_aw_bits_addr = axi4buf_1_auto_out_aw_bits_addr; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_aw_bits_len = axi4buf_1_auto_out_aw_bits_len; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_aw_bits_size = axi4buf_1_auto_out_aw_bits_size; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_aw_bits_burst = axi4buf_1_auto_out_aw_bits_burst; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_aw_bits_lock = axi4buf_1_auto_out_aw_bits_lock; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_aw_bits_cache = axi4buf_1_auto_out_aw_bits_cache; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_aw_bits_prot = axi4buf_1_auto_out_aw_bits_prot; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_aw_bits_qos = axi4buf_1_auto_out_aw_bits_qos; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_aw_bits_echo_tl_state_source = axi4buf_1_auto_out_aw_bits_echo_tl_state_source; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_w_valid = axi4buf_1_auto_out_w_valid; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_w_bits_data = axi4buf_1_auto_out_w_bits_data; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_w_bits_strb = axi4buf_1_auto_out_w_bits_strb; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_w_bits_last = axi4buf_1_auto_out_w_bits_last; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_b_ready = axi4buf_1_auto_out_b_ready; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_ar_valid = axi4buf_1_auto_out_ar_valid; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_ar_bits_id = axi4buf_1_auto_out_ar_bits_id; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_ar_bits_addr = axi4buf_1_auto_out_ar_bits_addr; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_ar_bits_len = axi4buf_1_auto_out_ar_bits_len; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_ar_bits_size = axi4buf_1_auto_out_ar_bits_size; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_ar_bits_burst = axi4buf_1_auto_out_ar_bits_burst; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_ar_bits_lock = axi4buf_1_auto_out_ar_bits_lock; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_ar_bits_cache = axi4buf_1_auto_out_ar_bits_cache; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_ar_bits_prot = axi4buf_1_auto_out_ar_bits_prot; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_ar_bits_qos = axi4buf_1_auto_out_ar_bits_qos; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_ar_bits_echo_tl_state_source = axi4buf_1_auto_out_ar_bits_echo_tl_state_source; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_in_r_ready = axi4buf_1_auto_out_r_ready; // @[LazyModule.scala 353:16]
  assign axi4buf_auto_out_aw_ready = axi4xbar_auto_in_0_aw_ready; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign axi4buf_auto_out_w_ready = axi4xbar_auto_in_0_w_ready; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign axi4buf_auto_out_b_valid = axi4xbar_auto_in_0_b_valid; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign axi4buf_auto_out_b_bits_id = axi4xbar_auto_in_0_b_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign axi4buf_auto_out_b_bits_echo_tl_state_source = axi4xbar_auto_in_0_b_bits_echo_tl_state_source; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign axi4buf_auto_out_ar_ready = axi4xbar_auto_in_0_ar_ready; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign axi4buf_auto_out_r_valid = axi4xbar_auto_in_0_r_valid; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign axi4buf_auto_out_r_bits_id = axi4xbar_auto_in_0_r_bits_id; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign axi4buf_auto_out_r_bits_data = axi4xbar_auto_in_0_r_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign axi4buf_auto_out_r_bits_echo_tl_state_source = axi4xbar_auto_in_0_r_bits_echo_tl_state_source; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign axi4buf_auto_out_r_bits_last = axi4xbar_auto_in_0_r_bits_last; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign axi4buf_1_clock = clock;
  assign axi4buf_1_reset = reset;
  assign axi4buf_1_auto_in_aw_valid = tl2axi4_auto_out_aw_valid; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_aw_bits_id = tl2axi4_auto_out_aw_bits_id; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_aw_bits_addr = tl2axi4_auto_out_aw_bits_addr; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_aw_bits_len = tl2axi4_auto_out_aw_bits_len; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_aw_bits_size = tl2axi4_auto_out_aw_bits_size; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_aw_bits_burst = tl2axi4_auto_out_aw_bits_burst; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_aw_bits_lock = tl2axi4_auto_out_aw_bits_lock; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_aw_bits_cache = tl2axi4_auto_out_aw_bits_cache; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_aw_bits_prot = tl2axi4_auto_out_aw_bits_prot; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_aw_bits_qos = tl2axi4_auto_out_aw_bits_qos; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_aw_bits_echo_tl_state_source = tl2axi4_auto_out_aw_bits_echo_tl_state_source; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_w_valid = tl2axi4_auto_out_w_valid; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_w_bits_data = tl2axi4_auto_out_w_bits_data; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_w_bits_strb = tl2axi4_auto_out_w_bits_strb; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_w_bits_last = tl2axi4_auto_out_w_bits_last; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_b_ready = tl2axi4_auto_out_b_ready; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_ar_valid = tl2axi4_auto_out_ar_valid; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_ar_bits_id = tl2axi4_auto_out_ar_bits_id; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_ar_bits_addr = tl2axi4_auto_out_ar_bits_addr; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_ar_bits_len = tl2axi4_auto_out_ar_bits_len; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_ar_bits_size = tl2axi4_auto_out_ar_bits_size; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_ar_bits_burst = tl2axi4_auto_out_ar_bits_burst; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_ar_bits_lock = tl2axi4_auto_out_ar_bits_lock; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_ar_bits_cache = tl2axi4_auto_out_ar_bits_cache; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_ar_bits_prot = tl2axi4_auto_out_ar_bits_prot; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_ar_bits_qos = tl2axi4_auto_out_ar_bits_qos; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_ar_bits_echo_tl_state_source = tl2axi4_auto_out_ar_bits_echo_tl_state_source; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_in_r_ready = tl2axi4_auto_out_r_ready; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_out_aw_ready = axi4buf_auto_in_aw_ready; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_out_w_ready = axi4buf_auto_in_w_ready; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_out_b_valid = axi4buf_auto_in_b_valid; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_out_b_bits_id = axi4buf_auto_in_b_bits_id; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_out_b_bits_echo_tl_state_source = axi4buf_auto_in_b_bits_echo_tl_state_source; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_out_ar_ready = axi4buf_auto_in_ar_ready; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_out_r_valid = axi4buf_auto_in_r_valid; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_out_r_bits_id = axi4buf_auto_in_r_bits_id; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_out_r_bits_data = axi4buf_auto_in_r_bits_data; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_out_r_bits_echo_tl_state_source = axi4buf_auto_in_r_bits_echo_tl_state_source; // @[LazyModule.scala 353:16]
  assign axi4buf_1_auto_out_r_bits_last = axi4buf_auto_in_r_bits_last; // @[LazyModule.scala 353:16]
  assign tl2axi4_clock = clock;
  assign tl2axi4_reset = reset;
  assign tl2axi4_auto_in_a_valid = acc_auto_mem_out_a_valid; // @[LazyModule.scala 355:16]
  assign tl2axi4_auto_in_a_bits_opcode = acc_auto_mem_out_a_bits_opcode; // @[LazyModule.scala 355:16]
  assign tl2axi4_auto_in_a_bits_size = acc_auto_mem_out_a_bits_size; // @[LazyModule.scala 355:16]
  assign tl2axi4_auto_in_a_bits_source = acc_auto_mem_out_a_bits_source; // @[LazyModule.scala 355:16]
  assign tl2axi4_auto_in_a_bits_address = acc_auto_mem_out_a_bits_address; // @[LazyModule.scala 355:16]
  assign tl2axi4_auto_in_a_bits_mask = acc_auto_mem_out_a_bits_mask; // @[LazyModule.scala 355:16]
  assign tl2axi4_auto_in_a_bits_data = acc_auto_mem_out_a_bits_data; // @[LazyModule.scala 355:16]
  assign tl2axi4_auto_in_d_ready = acc_auto_mem_out_d_ready; // @[LazyModule.scala 355:16]
  assign tl2axi4_auto_out_aw_ready = axi4buf_1_auto_in_aw_ready; // @[LazyModule.scala 353:16]
  assign tl2axi4_auto_out_w_ready = axi4buf_1_auto_in_w_ready; // @[LazyModule.scala 353:16]
  assign tl2axi4_auto_out_b_valid = axi4buf_1_auto_in_b_valid; // @[LazyModule.scala 353:16]
  assign tl2axi4_auto_out_b_bits_id = axi4buf_1_auto_in_b_bits_id; // @[LazyModule.scala 353:16]
  assign tl2axi4_auto_out_b_bits_echo_tl_state_source = axi4buf_1_auto_in_b_bits_echo_tl_state_source; // @[LazyModule.scala 353:16]
  assign tl2axi4_auto_out_ar_ready = axi4buf_1_auto_in_ar_ready; // @[LazyModule.scala 353:16]
  assign tl2axi4_auto_out_r_valid = axi4buf_1_auto_in_r_valid; // @[LazyModule.scala 353:16]
  assign tl2axi4_auto_out_r_bits_id = axi4buf_1_auto_in_r_bits_id; // @[LazyModule.scala 353:16]
  assign tl2axi4_auto_out_r_bits_data = axi4buf_1_auto_in_r_bits_data; // @[LazyModule.scala 353:16]
  assign tl2axi4_auto_out_r_bits_echo_tl_state_source = axi4buf_1_auto_in_r_bits_echo_tl_state_source; // @[LazyModule.scala 353:16]
  assign tl2axi4_auto_out_r_bits_last = axi4buf_1_auto_in_r_bits_last; // @[LazyModule.scala 353:16]
  assign axi4xbar_clock = clock;
  assign axi4xbar_reset = reset;
  assign axi4xbar_auto_in_1_aw_valid = axi4xbar_1_auto_out_aw_valid; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_aw_bits_id = axi4xbar_1_auto_out_aw_bits_id; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_aw_bits_addr = axi4xbar_1_auto_out_aw_bits_addr; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_aw_bits_len = axi4xbar_1_auto_out_aw_bits_len; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_aw_bits_size = axi4xbar_1_auto_out_aw_bits_size; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_aw_bits_burst = axi4xbar_1_auto_out_aw_bits_burst; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_aw_bits_lock = axi4xbar_1_auto_out_aw_bits_lock; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_aw_bits_cache = axi4xbar_1_auto_out_aw_bits_cache; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_aw_bits_prot = axi4xbar_1_auto_out_aw_bits_prot; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_aw_bits_qos = axi4xbar_1_auto_out_aw_bits_qos; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_w_valid = axi4xbar_1_auto_out_w_valid; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_w_bits_data = axi4xbar_1_auto_out_w_bits_data; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_w_bits_strb = axi4xbar_1_auto_out_w_bits_strb; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_w_bits_last = axi4xbar_1_auto_out_w_bits_last; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_b_ready = axi4xbar_1_auto_out_b_ready; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_ar_valid = axi4xbar_1_auto_out_ar_valid; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_ar_bits_id = axi4xbar_1_auto_out_ar_bits_id; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_ar_bits_addr = axi4xbar_1_auto_out_ar_bits_addr; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_ar_bits_len = axi4xbar_1_auto_out_ar_bits_len; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_ar_bits_size = axi4xbar_1_auto_out_ar_bits_size; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_ar_bits_burst = axi4xbar_1_auto_out_ar_bits_burst; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_ar_bits_lock = axi4xbar_1_auto_out_ar_bits_lock; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_ar_bits_cache = axi4xbar_1_auto_out_ar_bits_cache; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_ar_bits_prot = axi4xbar_1_auto_out_ar_bits_prot; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_ar_bits_qos = axi4xbar_1_auto_out_ar_bits_qos; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_1_r_ready = axi4xbar_1_auto_out_r_ready; // @[LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_aw_valid = axi4buf_auto_out_aw_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_aw_bits_id = axi4buf_auto_out_aw_bits_id; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_aw_bits_addr = axi4buf_auto_out_aw_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_aw_bits_len = axi4buf_auto_out_aw_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_aw_bits_size = axi4buf_auto_out_aw_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_aw_bits_burst = axi4buf_auto_out_aw_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_aw_bits_lock = axi4buf_auto_out_aw_bits_lock; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_aw_bits_cache = axi4buf_auto_out_aw_bits_cache; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_aw_bits_prot = axi4buf_auto_out_aw_bits_prot; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_aw_bits_qos = axi4buf_auto_out_aw_bits_qos; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_aw_bits_echo_tl_state_source = axi4buf_auto_out_aw_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_w_valid = axi4buf_auto_out_w_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_w_bits_data = axi4buf_auto_out_w_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_w_bits_strb = axi4buf_auto_out_w_bits_strb; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_w_bits_last = axi4buf_auto_out_w_bits_last; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_b_ready = axi4buf_auto_out_b_ready; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_ar_valid = axi4buf_auto_out_ar_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_ar_bits_id = axi4buf_auto_out_ar_bits_id; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_ar_bits_addr = axi4buf_auto_out_ar_bits_addr; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_ar_bits_len = axi4buf_auto_out_ar_bits_len; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_ar_bits_size = axi4buf_auto_out_ar_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_ar_bits_burst = axi4buf_auto_out_ar_bits_burst; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_ar_bits_lock = axi4buf_auto_out_ar_bits_lock; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_ar_bits_cache = axi4buf_auto_out_ar_bits_cache; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_ar_bits_prot = axi4buf_auto_out_ar_bits_prot; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_ar_bits_qos = axi4buf_auto_out_ar_bits_qos; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_ar_bits_echo_tl_state_source = axi4buf_auto_out_ar_bits_echo_tl_state_source; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_in_0_r_ready = axi4buf_auto_out_r_ready; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign axi4xbar_auto_out_aw_ready = axi4buf_5_auto_in_aw_ready; // @[LazyModule.scala 355:16]
  assign axi4xbar_auto_out_w_ready = axi4buf_5_auto_in_w_ready; // @[LazyModule.scala 355:16]
  assign axi4xbar_auto_out_b_valid = axi4buf_5_auto_in_b_valid; // @[LazyModule.scala 355:16]
  assign axi4xbar_auto_out_b_bits_id = axi4buf_5_auto_in_b_bits_id; // @[LazyModule.scala 355:16]
  assign axi4xbar_auto_out_b_bits_resp = axi4buf_5_auto_in_b_bits_resp; // @[LazyModule.scala 355:16]
  assign axi4xbar_auto_out_b_bits_echo_tl_state_source = axi4buf_5_auto_in_b_bits_echo_tl_state_source; // @[LazyModule.scala 355:16]
  assign axi4xbar_auto_out_ar_ready = axi4buf_5_auto_in_ar_ready; // @[LazyModule.scala 355:16]
  assign axi4xbar_auto_out_r_valid = axi4buf_5_auto_in_r_valid; // @[LazyModule.scala 355:16]
  assign axi4xbar_auto_out_r_bits_id = axi4buf_5_auto_in_r_bits_id; // @[LazyModule.scala 355:16]
  assign axi4xbar_auto_out_r_bits_data = axi4buf_5_auto_in_r_bits_data; // @[LazyModule.scala 355:16]
  assign axi4xbar_auto_out_r_bits_resp = axi4buf_5_auto_in_r_bits_resp; // @[LazyModule.scala 355:16]
  assign axi4xbar_auto_out_r_bits_echo_tl_state_source = axi4buf_5_auto_in_r_bits_echo_tl_state_source; // @[LazyModule.scala 355:16]
  assign axi4xbar_auto_out_r_bits_last = axi4buf_5_auto_in_r_bits_last; // @[LazyModule.scala 355:16]
  assign axi4xbar_1_clock = clock;
  assign axi4xbar_1_reset = reset;
  assign axi4xbar_1_auto_in_aw_valid = axi4buf_2_auto_out_aw_valid; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_aw_bits_id = axi4buf_2_auto_out_aw_bits_id; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_aw_bits_addr = axi4buf_2_auto_out_aw_bits_addr; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_aw_bits_len = axi4buf_2_auto_out_aw_bits_len; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_aw_bits_size = axi4buf_2_auto_out_aw_bits_size; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_aw_bits_burst = axi4buf_2_auto_out_aw_bits_burst; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_aw_bits_lock = axi4buf_2_auto_out_aw_bits_lock; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_aw_bits_cache = axi4buf_2_auto_out_aw_bits_cache; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_aw_bits_prot = axi4buf_2_auto_out_aw_bits_prot; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_aw_bits_qos = axi4buf_2_auto_out_aw_bits_qos; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_w_valid = axi4buf_2_auto_out_w_valid; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_w_bits_data = axi4buf_2_auto_out_w_bits_data; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_w_bits_strb = axi4buf_2_auto_out_w_bits_strb; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_w_bits_last = axi4buf_2_auto_out_w_bits_last; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_b_ready = axi4buf_2_auto_out_b_ready; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_ar_valid = axi4buf_2_auto_out_ar_valid; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_ar_bits_id = axi4buf_2_auto_out_ar_bits_id; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_ar_bits_addr = axi4buf_2_auto_out_ar_bits_addr; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_ar_bits_len = axi4buf_2_auto_out_ar_bits_len; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_ar_bits_size = axi4buf_2_auto_out_ar_bits_size; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_ar_bits_burst = axi4buf_2_auto_out_ar_bits_burst; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_ar_bits_lock = axi4buf_2_auto_out_ar_bits_lock; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_ar_bits_cache = axi4buf_2_auto_out_ar_bits_cache; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_ar_bits_prot = axi4buf_2_auto_out_ar_bits_prot; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_ar_bits_qos = axi4buf_2_auto_out_ar_bits_qos; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_in_r_ready = axi4buf_2_auto_out_r_ready; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_out_aw_ready = axi4xbar_auto_in_1_aw_ready; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_out_w_ready = axi4xbar_auto_in_1_w_ready; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_out_b_valid = axi4xbar_auto_in_1_b_valid; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_out_b_bits_id = axi4xbar_auto_in_1_b_bits_id; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_out_b_bits_resp = axi4xbar_auto_in_1_b_bits_resp; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_out_ar_ready = axi4xbar_auto_in_1_ar_ready; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_out_r_valid = axi4xbar_auto_in_1_r_valid; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_out_r_bits_id = axi4xbar_auto_in_1_r_bits_id; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_out_r_bits_data = axi4xbar_auto_in_1_r_bits_data; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_out_r_bits_resp = axi4xbar_auto_in_1_r_bits_resp; // @[LazyModule.scala 353:16]
  assign axi4xbar_1_auto_out_r_bits_last = axi4xbar_auto_in_1_r_bits_last; // @[LazyModule.scala 353:16]
  assign axi4buf_2_clock = clock;
  assign axi4buf_2_reset = reset;
  assign axi4buf_2_auto_in_aw_valid = dma_awvalid; // @[Nodes.scala 1212:84 AXI4Compat.scala 131:19]
  assign axi4buf_2_auto_in_aw_bits_id = dma_awid; // @[AXI4Compat.scala 121:21 Nodes.scala 1212:84]
  assign axi4buf_2_auto_in_aw_bits_addr = dma_awaddr; // @[Nodes.scala 1212:84 AXI4Compat.scala 126:23]
  assign axi4buf_2_auto_in_aw_bits_len = dma_awlen; // @[Nodes.scala 1212:84 AXI4Compat.scala 123:22]
  assign axi4buf_2_auto_in_aw_bits_size = dma_awsize; // @[Nodes.scala 1212:84 AXI4Compat.scala 129:23]
  assign axi4buf_2_auto_in_aw_bits_burst = dma_awburst; // @[Nodes.scala 1212:84 AXI4Compat.scala 127:24]
  assign axi4buf_2_auto_in_aw_bits_lock = dma_awlock; // @[Nodes.scala 1212:84 AXI4Compat.scala 124:23]
  assign axi4buf_2_auto_in_aw_bits_cache = dma_awcache; // @[Nodes.scala 1212:84 AXI4Compat.scala 128:24]
  assign axi4buf_2_auto_in_aw_bits_prot = dma_awprot; // @[Nodes.scala 1212:84 AXI4Compat.scala 125:23]
  assign axi4buf_2_auto_in_aw_bits_qos = dma_awqos; // @[Nodes.scala 1212:84 AXI4Compat.scala 122:22]
  assign axi4buf_2_auto_in_w_valid = dma_wvalid; // @[Nodes.scala 1212:84 AXI4Compat.scala 141:18]
  assign axi4buf_2_auto_in_w_bits_data = dma_wdata; // @[Nodes.scala 1212:84 AXI4Compat.scala 138:22]
  assign axi4buf_2_auto_in_w_bits_strb = dma_wstrb; // @[Nodes.scala 1212:84 AXI4Compat.scala 139:22]
  assign axi4buf_2_auto_in_w_bits_last = dma_wlast; // @[Nodes.scala 1212:84 AXI4Compat.scala 140:22]
  assign axi4buf_2_auto_in_b_ready = dma_bready; // @[Nodes.scala 1212:84 AXI4Compat.scala 135:18]
  assign axi4buf_2_auto_in_ar_valid = dma_arvalid; // @[AXI4Compat.scala 119:19 Nodes.scala 1212:84]
  assign axi4buf_2_auto_in_ar_bits_id = dma_arid; // @[AXI4Compat.scala 109:21 Nodes.scala 1212:84]
  assign axi4buf_2_auto_in_ar_bits_addr = dma_araddr; // @[AXI4Compat.scala 114:23 Nodes.scala 1212:84]
  assign axi4buf_2_auto_in_ar_bits_len = dma_arlen; // @[AXI4Compat.scala 111:22 Nodes.scala 1212:84]
  assign axi4buf_2_auto_in_ar_bits_size = dma_arsize; // @[AXI4Compat.scala 117:23 Nodes.scala 1212:84]
  assign axi4buf_2_auto_in_ar_bits_burst = dma_arburst; // @[AXI4Compat.scala 115:24 Nodes.scala 1212:84]
  assign axi4buf_2_auto_in_ar_bits_lock = dma_arlock; // @[AXI4Compat.scala 112:23 Nodes.scala 1212:84]
  assign axi4buf_2_auto_in_ar_bits_cache = dma_arcache; // @[AXI4Compat.scala 116:24 Nodes.scala 1212:84]
  assign axi4buf_2_auto_in_ar_bits_prot = dma_arprot; // @[AXI4Compat.scala 113:23 Nodes.scala 1212:84]
  assign axi4buf_2_auto_in_ar_bits_qos = dma_arqos; // @[AXI4Compat.scala 110:22 Nodes.scala 1212:84]
  assign axi4buf_2_auto_in_r_ready = dma_rready; // @[AXI4Compat.scala 107:18 Nodes.scala 1212:84]
  assign axi4buf_2_auto_out_aw_ready = axi4xbar_1_auto_in_aw_ready; // @[LazyModule.scala 353:16]
  assign axi4buf_2_auto_out_w_ready = axi4xbar_1_auto_in_w_ready; // @[LazyModule.scala 353:16]
  assign axi4buf_2_auto_out_b_valid = axi4xbar_1_auto_in_b_valid; // @[LazyModule.scala 353:16]
  assign axi4buf_2_auto_out_b_bits_id = axi4xbar_1_auto_in_b_bits_id; // @[LazyModule.scala 353:16]
  assign axi4buf_2_auto_out_b_bits_resp = axi4xbar_1_auto_in_b_bits_resp; // @[LazyModule.scala 353:16]
  assign axi4buf_2_auto_out_ar_ready = axi4xbar_1_auto_in_ar_ready; // @[LazyModule.scala 353:16]
  assign axi4buf_2_auto_out_r_valid = axi4xbar_1_auto_in_r_valid; // @[LazyModule.scala 353:16]
  assign axi4buf_2_auto_out_r_bits_id = axi4xbar_1_auto_in_r_bits_id; // @[LazyModule.scala 353:16]
  assign axi4buf_2_auto_out_r_bits_data = axi4xbar_1_auto_in_r_bits_data; // @[LazyModule.scala 353:16]
  assign axi4buf_2_auto_out_r_bits_resp = axi4xbar_1_auto_in_r_bits_resp; // @[LazyModule.scala 353:16]
  assign axi4buf_2_auto_out_r_bits_last = axi4xbar_1_auto_in_r_bits_last; // @[LazyModule.scala 353:16]
  assign axi4buf_3_clock = clock;
  assign axi4buf_3_reset = reset;
  assign axi4buf_3_auto_in_aw_valid = axi4yank_auto_out_aw_valid; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_aw_bits_id = axi4yank_auto_out_aw_bits_id; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_aw_bits_addr = axi4yank_auto_out_aw_bits_addr; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_aw_bits_len = axi4yank_auto_out_aw_bits_len; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_aw_bits_size = axi4yank_auto_out_aw_bits_size; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_aw_bits_burst = axi4yank_auto_out_aw_bits_burst; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_aw_bits_lock = axi4yank_auto_out_aw_bits_lock; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_aw_bits_cache = axi4yank_auto_out_aw_bits_cache; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_aw_bits_prot = axi4yank_auto_out_aw_bits_prot; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_aw_bits_qos = axi4yank_auto_out_aw_bits_qos; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_w_valid = axi4yank_auto_out_w_valid; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_w_bits_data = axi4yank_auto_out_w_bits_data; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_w_bits_strb = axi4yank_auto_out_w_bits_strb; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_w_bits_last = axi4yank_auto_out_w_bits_last; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_b_ready = axi4yank_auto_out_b_ready; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_ar_valid = axi4yank_auto_out_ar_valid; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_ar_bits_id = axi4yank_auto_out_ar_bits_id; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_ar_bits_addr = axi4yank_auto_out_ar_bits_addr; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_ar_bits_len = axi4yank_auto_out_ar_bits_len; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_ar_bits_size = axi4yank_auto_out_ar_bits_size; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_ar_bits_burst = axi4yank_auto_out_ar_bits_burst; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_ar_bits_lock = axi4yank_auto_out_ar_bits_lock; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_ar_bits_cache = axi4yank_auto_out_ar_bits_cache; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_ar_bits_prot = axi4yank_auto_out_ar_bits_prot; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_ar_bits_qos = axi4yank_auto_out_ar_bits_qos; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_in_r_ready = axi4yank_auto_out_r_ready; // @[LazyModule.scala 353:16]
  assign axi4buf_3_auto_out_aw_ready = M00_AXI_awready; // @[Nodes.scala 1215:84 AXI4Compat.scala 91:19]
  assign axi4buf_3_auto_out_w_ready = M00_AXI_wready; // @[Nodes.scala 1215:84 AXI4Compat.scala 98:18]
  assign axi4buf_3_auto_out_b_valid = M00_AXI_bvalid; // @[Nodes.scala 1215:84 AXI4Compat.scala 79:18]
  assign axi4buf_3_auto_out_b_bits_id = M00_AXI_bid; // @[Nodes.scala 1215:84 AXI4Compat.scala 76:20]
  assign axi4buf_3_auto_out_b_bits_resp = M00_AXI_bresp; // @[Nodes.scala 1215:84 AXI4Compat.scala 77:22]
  assign axi4buf_3_auto_out_ar_ready = M00_AXI_arready; // @[Nodes.scala 1215:84 AXI4Compat.scala 73:19]
  assign axi4buf_3_auto_out_r_valid = M00_AXI_rvalid; // @[Nodes.scala 1215:84 AXI4Compat.scala 60:18]
  assign axi4buf_3_auto_out_r_bits_id = M00_AXI_rid; // @[Nodes.scala 1215:84 AXI4Compat.scala 56:20]
  assign axi4buf_3_auto_out_r_bits_data = M00_AXI_rdata; // @[Nodes.scala 1215:84 AXI4Compat.scala 57:22]
  assign axi4buf_3_auto_out_r_bits_resp = M00_AXI_rresp; // @[Nodes.scala 1215:84 AXI4Compat.scala 58:22]
  assign axi4buf_3_auto_out_r_bits_last = M00_AXI_rlast; // @[Nodes.scala 1215:84 AXI4Compat.scala 59:22]
  assign axi4yank_clock = clock;
  assign axi4yank_reset = reset;
  assign axi4yank_auto_in_aw_valid = axi4buf_4_auto_out_aw_valid; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_aw_bits_id = axi4buf_4_auto_out_aw_bits_id; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_aw_bits_addr = axi4buf_4_auto_out_aw_bits_addr; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_aw_bits_len = axi4buf_4_auto_out_aw_bits_len; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_aw_bits_size = axi4buf_4_auto_out_aw_bits_size; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_aw_bits_burst = axi4buf_4_auto_out_aw_bits_burst; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_aw_bits_lock = axi4buf_4_auto_out_aw_bits_lock; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_aw_bits_cache = axi4buf_4_auto_out_aw_bits_cache; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_aw_bits_prot = axi4buf_4_auto_out_aw_bits_prot; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_aw_bits_qos = axi4buf_4_auto_out_aw_bits_qos; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_aw_bits_echo_tl_state_source = axi4buf_4_auto_out_aw_bits_echo_tl_state_source; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_aw_bits_echo_extra_id = axi4buf_4_auto_out_aw_bits_echo_extra_id; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_w_valid = axi4buf_4_auto_out_w_valid; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_w_bits_data = axi4buf_4_auto_out_w_bits_data; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_w_bits_strb = axi4buf_4_auto_out_w_bits_strb; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_w_bits_last = axi4buf_4_auto_out_w_bits_last; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_b_ready = axi4buf_4_auto_out_b_ready; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_ar_valid = axi4buf_4_auto_out_ar_valid; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_ar_bits_id = axi4buf_4_auto_out_ar_bits_id; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_ar_bits_addr = axi4buf_4_auto_out_ar_bits_addr; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_ar_bits_len = axi4buf_4_auto_out_ar_bits_len; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_ar_bits_size = axi4buf_4_auto_out_ar_bits_size; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_ar_bits_burst = axi4buf_4_auto_out_ar_bits_burst; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_ar_bits_lock = axi4buf_4_auto_out_ar_bits_lock; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_ar_bits_cache = axi4buf_4_auto_out_ar_bits_cache; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_ar_bits_prot = axi4buf_4_auto_out_ar_bits_prot; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_ar_bits_qos = axi4buf_4_auto_out_ar_bits_qos; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_ar_bits_echo_tl_state_source = axi4buf_4_auto_out_ar_bits_echo_tl_state_source; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_ar_bits_echo_extra_id = axi4buf_4_auto_out_ar_bits_echo_extra_id; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_in_r_ready = axi4buf_4_auto_out_r_ready; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_out_aw_ready = axi4buf_3_auto_in_aw_ready; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_out_w_ready = axi4buf_3_auto_in_w_ready; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_out_b_valid = axi4buf_3_auto_in_b_valid; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_out_b_bits_id = axi4buf_3_auto_in_b_bits_id; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_out_b_bits_resp = axi4buf_3_auto_in_b_bits_resp; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_out_ar_ready = axi4buf_3_auto_in_ar_ready; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_out_r_valid = axi4buf_3_auto_in_r_valid; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_out_r_bits_id = axi4buf_3_auto_in_r_bits_id; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_out_r_bits_data = axi4buf_3_auto_in_r_bits_data; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_out_r_bits_resp = axi4buf_3_auto_in_r_bits_resp; // @[LazyModule.scala 353:16]
  assign axi4yank_auto_out_r_bits_last = axi4buf_3_auto_in_r_bits_last; // @[LazyModule.scala 353:16]
  assign axi4buf_4_clock = clock;
  assign axi4buf_4_reset = reset;
  assign axi4buf_4_auto_in_aw_valid = axi4index_auto_out_aw_valid; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_aw_bits_id = axi4index_auto_out_aw_bits_id; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_aw_bits_addr = axi4index_auto_out_aw_bits_addr; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_aw_bits_len = axi4index_auto_out_aw_bits_len; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_aw_bits_size = axi4index_auto_out_aw_bits_size; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_aw_bits_burst = axi4index_auto_out_aw_bits_burst; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_aw_bits_lock = axi4index_auto_out_aw_bits_lock; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_aw_bits_cache = axi4index_auto_out_aw_bits_cache; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_aw_bits_prot = axi4index_auto_out_aw_bits_prot; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_aw_bits_qos = axi4index_auto_out_aw_bits_qos; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_aw_bits_echo_tl_state_source = axi4index_auto_out_aw_bits_echo_tl_state_source; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_aw_bits_echo_extra_id = axi4index_auto_out_aw_bits_echo_extra_id; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_w_valid = axi4index_auto_out_w_valid; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_w_bits_data = axi4index_auto_out_w_bits_data; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_w_bits_strb = axi4index_auto_out_w_bits_strb; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_w_bits_last = axi4index_auto_out_w_bits_last; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_b_ready = axi4index_auto_out_b_ready; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_ar_valid = axi4index_auto_out_ar_valid; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_ar_bits_id = axi4index_auto_out_ar_bits_id; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_ar_bits_addr = axi4index_auto_out_ar_bits_addr; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_ar_bits_len = axi4index_auto_out_ar_bits_len; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_ar_bits_size = axi4index_auto_out_ar_bits_size; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_ar_bits_burst = axi4index_auto_out_ar_bits_burst; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_ar_bits_lock = axi4index_auto_out_ar_bits_lock; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_ar_bits_cache = axi4index_auto_out_ar_bits_cache; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_ar_bits_prot = axi4index_auto_out_ar_bits_prot; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_ar_bits_qos = axi4index_auto_out_ar_bits_qos; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_ar_bits_echo_tl_state_source = axi4index_auto_out_ar_bits_echo_tl_state_source; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_ar_bits_echo_extra_id = axi4index_auto_out_ar_bits_echo_extra_id; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_in_r_ready = axi4index_auto_out_r_ready; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_out_aw_ready = axi4yank_auto_in_aw_ready; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_out_w_ready = axi4yank_auto_in_w_ready; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_out_b_valid = axi4yank_auto_in_b_valid; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_out_b_bits_id = axi4yank_auto_in_b_bits_id; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_out_b_bits_resp = axi4yank_auto_in_b_bits_resp; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_out_b_bits_echo_tl_state_source = axi4yank_auto_in_b_bits_echo_tl_state_source; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_out_b_bits_echo_extra_id = axi4yank_auto_in_b_bits_echo_extra_id; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_out_ar_ready = axi4yank_auto_in_ar_ready; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_out_r_valid = axi4yank_auto_in_r_valid; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_out_r_bits_id = axi4yank_auto_in_r_bits_id; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_out_r_bits_data = axi4yank_auto_in_r_bits_data; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_out_r_bits_resp = axi4yank_auto_in_r_bits_resp; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_out_r_bits_echo_tl_state_source = axi4yank_auto_in_r_bits_echo_tl_state_source; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_out_r_bits_echo_extra_id = axi4yank_auto_in_r_bits_echo_extra_id; // @[LazyModule.scala 353:16]
  assign axi4buf_4_auto_out_r_bits_last = axi4yank_auto_in_r_bits_last; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_aw_valid = axi4buf_5_auto_out_aw_valid; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_aw_bits_id = axi4buf_5_auto_out_aw_bits_id; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_aw_bits_addr = axi4buf_5_auto_out_aw_bits_addr; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_aw_bits_len = axi4buf_5_auto_out_aw_bits_len; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_aw_bits_size = axi4buf_5_auto_out_aw_bits_size; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_aw_bits_burst = axi4buf_5_auto_out_aw_bits_burst; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_aw_bits_lock = axi4buf_5_auto_out_aw_bits_lock; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_aw_bits_cache = axi4buf_5_auto_out_aw_bits_cache; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_aw_bits_prot = axi4buf_5_auto_out_aw_bits_prot; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_aw_bits_qos = axi4buf_5_auto_out_aw_bits_qos; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_aw_bits_echo_tl_state_source = axi4buf_5_auto_out_aw_bits_echo_tl_state_source; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_w_valid = axi4buf_5_auto_out_w_valid; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_w_bits_data = axi4buf_5_auto_out_w_bits_data; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_w_bits_strb = axi4buf_5_auto_out_w_bits_strb; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_w_bits_last = axi4buf_5_auto_out_w_bits_last; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_b_ready = axi4buf_5_auto_out_b_ready; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_ar_valid = axi4buf_5_auto_out_ar_valid; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_ar_bits_id = axi4buf_5_auto_out_ar_bits_id; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_ar_bits_addr = axi4buf_5_auto_out_ar_bits_addr; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_ar_bits_len = axi4buf_5_auto_out_ar_bits_len; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_ar_bits_size = axi4buf_5_auto_out_ar_bits_size; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_ar_bits_burst = axi4buf_5_auto_out_ar_bits_burst; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_ar_bits_lock = axi4buf_5_auto_out_ar_bits_lock; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_ar_bits_cache = axi4buf_5_auto_out_ar_bits_cache; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_ar_bits_prot = axi4buf_5_auto_out_ar_bits_prot; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_ar_bits_qos = axi4buf_5_auto_out_ar_bits_qos; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_ar_bits_echo_tl_state_source = axi4buf_5_auto_out_ar_bits_echo_tl_state_source; // @[LazyModule.scala 353:16]
  assign axi4index_auto_in_r_ready = axi4buf_5_auto_out_r_ready; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_aw_ready = axi4buf_4_auto_in_aw_ready; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_w_ready = axi4buf_4_auto_in_w_ready; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_b_valid = axi4buf_4_auto_in_b_valid; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_b_bits_id = axi4buf_4_auto_in_b_bits_id; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_b_bits_resp = axi4buf_4_auto_in_b_bits_resp; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_b_bits_echo_tl_state_source = axi4buf_4_auto_in_b_bits_echo_tl_state_source; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_b_bits_echo_extra_id = axi4buf_4_auto_in_b_bits_echo_extra_id; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_ar_ready = axi4buf_4_auto_in_ar_ready; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_r_valid = axi4buf_4_auto_in_r_valid; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_r_bits_id = axi4buf_4_auto_in_r_bits_id; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_r_bits_data = axi4buf_4_auto_in_r_bits_data; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_r_bits_resp = axi4buf_4_auto_in_r_bits_resp; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_r_bits_echo_tl_state_source = axi4buf_4_auto_in_r_bits_echo_tl_state_source; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_r_bits_echo_extra_id = axi4buf_4_auto_in_r_bits_echo_extra_id; // @[LazyModule.scala 353:16]
  assign axi4index_auto_out_r_bits_last = axi4buf_4_auto_in_r_bits_last; // @[LazyModule.scala 353:16]
  assign axi4buf_5_clock = clock;
  assign axi4buf_5_reset = reset;
  assign axi4buf_5_auto_in_aw_valid = axi4xbar_auto_out_aw_valid; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_aw_bits_id = axi4xbar_auto_out_aw_bits_id; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_aw_bits_addr = axi4xbar_auto_out_aw_bits_addr; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_aw_bits_len = axi4xbar_auto_out_aw_bits_len; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_aw_bits_size = axi4xbar_auto_out_aw_bits_size; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_aw_bits_burst = axi4xbar_auto_out_aw_bits_burst; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_aw_bits_lock = axi4xbar_auto_out_aw_bits_lock; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_aw_bits_cache = axi4xbar_auto_out_aw_bits_cache; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_aw_bits_prot = axi4xbar_auto_out_aw_bits_prot; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_aw_bits_qos = axi4xbar_auto_out_aw_bits_qos; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_aw_bits_echo_tl_state_source = axi4xbar_auto_out_aw_bits_echo_tl_state_source; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_w_valid = axi4xbar_auto_out_w_valid; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_w_bits_data = axi4xbar_auto_out_w_bits_data; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_w_bits_strb = axi4xbar_auto_out_w_bits_strb; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_w_bits_last = axi4xbar_auto_out_w_bits_last; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_b_ready = axi4xbar_auto_out_b_ready; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_ar_valid = axi4xbar_auto_out_ar_valid; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_ar_bits_id = axi4xbar_auto_out_ar_bits_id; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_ar_bits_addr = axi4xbar_auto_out_ar_bits_addr; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_ar_bits_len = axi4xbar_auto_out_ar_bits_len; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_ar_bits_size = axi4xbar_auto_out_ar_bits_size; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_ar_bits_burst = axi4xbar_auto_out_ar_bits_burst; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_ar_bits_lock = axi4xbar_auto_out_ar_bits_lock; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_ar_bits_cache = axi4xbar_auto_out_ar_bits_cache; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_ar_bits_prot = axi4xbar_auto_out_ar_bits_prot; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_ar_bits_qos = axi4xbar_auto_out_ar_bits_qos; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_ar_bits_echo_tl_state_source = axi4xbar_auto_out_ar_bits_echo_tl_state_source; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_in_r_ready = axi4xbar_auto_out_r_ready; // @[LazyModule.scala 355:16]
  assign axi4buf_5_auto_out_aw_ready = axi4index_auto_in_aw_ready; // @[LazyModule.scala 353:16]
  assign axi4buf_5_auto_out_w_ready = axi4index_auto_in_w_ready; // @[LazyModule.scala 353:16]
  assign axi4buf_5_auto_out_b_valid = axi4index_auto_in_b_valid; // @[LazyModule.scala 353:16]
  assign axi4buf_5_auto_out_b_bits_id = axi4index_auto_in_b_bits_id; // @[LazyModule.scala 353:16]
  assign axi4buf_5_auto_out_b_bits_resp = axi4index_auto_in_b_bits_resp; // @[LazyModule.scala 353:16]
  assign axi4buf_5_auto_out_b_bits_echo_tl_state_source = axi4index_auto_in_b_bits_echo_tl_state_source; // @[LazyModule.scala 353:16]
  assign axi4buf_5_auto_out_ar_ready = axi4index_auto_in_ar_ready; // @[LazyModule.scala 353:16]
  assign axi4buf_5_auto_out_r_valid = axi4index_auto_in_r_valid; // @[LazyModule.scala 353:16]
  assign axi4buf_5_auto_out_r_bits_id = axi4index_auto_in_r_bits_id; // @[LazyModule.scala 353:16]
  assign axi4buf_5_auto_out_r_bits_data = axi4index_auto_in_r_bits_data; // @[LazyModule.scala 353:16]
  assign axi4buf_5_auto_out_r_bits_resp = axi4index_auto_in_r_bits_resp; // @[LazyModule.scala 353:16]
  assign axi4buf_5_auto_out_r_bits_echo_tl_state_source = axi4index_auto_in_r_bits_echo_tl_state_source; // @[LazyModule.scala 353:16]
  assign axi4buf_5_auto_out_r_bits_last = axi4index_auto_in_r_bits_last; // @[LazyModule.scala 353:16]
  assign cmd_resp_axilhub_clock = clock;
  assign cmd_resp_axilhub_reset = reset;
  assign cmd_resp_axilhub_auto_in_aw_valid = axi4buf_6_auto_out_aw_valid; // @[LazyModule.scala 353:16]
  assign cmd_resp_axilhub_auto_in_aw_bits_id = axi4buf_6_auto_out_aw_bits_id; // @[LazyModule.scala 353:16]
  assign cmd_resp_axilhub_auto_in_aw_bits_addr = axi4buf_6_auto_out_aw_bits_addr; // @[LazyModule.scala 353:16]
  assign cmd_resp_axilhub_auto_in_aw_bits_len = axi4buf_6_auto_out_aw_bits_len; // @[LazyModule.scala 353:16]
  assign cmd_resp_axilhub_auto_in_aw_bits_size = axi4buf_6_auto_out_aw_bits_size; // @[LazyModule.scala 353:16]
  assign cmd_resp_axilhub_auto_in_aw_bits_burst = axi4buf_6_auto_out_aw_bits_burst; // @[LazyModule.scala 353:16]
  assign cmd_resp_axilhub_auto_in_w_valid = axi4buf_6_auto_out_w_valid; // @[LazyModule.scala 353:16]
  assign cmd_resp_axilhub_auto_in_w_bits_data = axi4buf_6_auto_out_w_bits_data; // @[LazyModule.scala 353:16]
  assign cmd_resp_axilhub_auto_in_w_bits_last = axi4buf_6_auto_out_w_bits_last; // @[LazyModule.scala 353:16]
  assign cmd_resp_axilhub_auto_in_b_ready = axi4buf_6_auto_out_b_ready; // @[LazyModule.scala 353:16]
  assign cmd_resp_axilhub_auto_in_ar_valid = axi4buf_6_auto_out_ar_valid; // @[LazyModule.scala 353:16]
  assign cmd_resp_axilhub_auto_in_ar_bits_id = axi4buf_6_auto_out_ar_bits_id; // @[LazyModule.scala 353:16]
  assign cmd_resp_axilhub_auto_in_ar_bits_addr = axi4buf_6_auto_out_ar_bits_addr; // @[LazyModule.scala 353:16]
  assign cmd_resp_axilhub_auto_in_ar_bits_len = axi4buf_6_auto_out_ar_bits_len; // @[LazyModule.scala 353:16]
  assign cmd_resp_axilhub_auto_in_ar_bits_size = axi4buf_6_auto_out_ar_bits_size; // @[LazyModule.scala 353:16]
  assign cmd_resp_axilhub_auto_in_ar_bits_burst = axi4buf_6_auto_out_ar_bits_burst; // @[LazyModule.scala 353:16]
  assign cmd_resp_axilhub_auto_in_r_ready = axi4buf_6_auto_out_r_ready; // @[LazyModule.scala 353:16]
  assign cmd_resp_axilhub_io_rocc_in_ready = acc_io_cmd_ready; // @[ComposerTop.scala 148:21]
  assign cmd_resp_axilhub_io_rocc_out_valid = acc_io_resp_valid; // @[ComposerTop.scala 149:31]
  assign cmd_resp_axilhub_io_rocc_out_bits_rd = acc_io_resp_bits_rd; // @[ComposerTop.scala 149:31]
  assign cmd_resp_axilhub_io_rocc_out_bits_data = 5'h10 == acc_io_resp_bits_rd ? arCnt : _GEN_12; // @[ComposerTop.scala 204:38 206:45]
  assign axi4buf_6_clock = clock;
  assign axi4buf_6_reset = reset;
  assign axi4buf_6_auto_in_aw_valid = S00_AXI_awvalid; // @[Nodes.scala 1212:84 AXI4Compat.scala 131:19]
  assign axi4buf_6_auto_in_aw_bits_id = S00_AXI_awid; // @[AXI4Compat.scala 121:21 Nodes.scala 1212:84]
  assign axi4buf_6_auto_in_aw_bits_addr = S00_AXI_awaddr; // @[Nodes.scala 1212:84 AXI4Compat.scala 126:23]
  assign axi4buf_6_auto_in_aw_bits_len = S00_AXI_awlen; // @[Nodes.scala 1212:84 AXI4Compat.scala 123:22]
  assign axi4buf_6_auto_in_aw_bits_size = S00_AXI_awsize; // @[Nodes.scala 1212:84 AXI4Compat.scala 129:23]
  assign axi4buf_6_auto_in_aw_bits_burst = S00_AXI_awburst; // @[Nodes.scala 1212:84 AXI4Compat.scala 127:24]
  assign axi4buf_6_auto_in_w_valid = S00_AXI_wvalid; // @[Nodes.scala 1212:84 AXI4Compat.scala 141:18]
  assign axi4buf_6_auto_in_w_bits_data = S00_AXI_wdata; // @[Nodes.scala 1212:84 AXI4Compat.scala 138:22]
  assign axi4buf_6_auto_in_w_bits_last = S00_AXI_wlast; // @[Nodes.scala 1212:84 AXI4Compat.scala 140:22]
  assign axi4buf_6_auto_in_b_ready = S00_AXI_bready; // @[Nodes.scala 1212:84 AXI4Compat.scala 135:18]
  assign axi4buf_6_auto_in_ar_valid = S00_AXI_arvalid; // @[AXI4Compat.scala 119:19 Nodes.scala 1212:84]
  assign axi4buf_6_auto_in_ar_bits_id = S00_AXI_arid; // @[AXI4Compat.scala 109:21 Nodes.scala 1212:84]
  assign axi4buf_6_auto_in_ar_bits_addr = S00_AXI_araddr; // @[AXI4Compat.scala 114:23 Nodes.scala 1212:84]
  assign axi4buf_6_auto_in_ar_bits_len = S00_AXI_arlen; // @[AXI4Compat.scala 111:22 Nodes.scala 1212:84]
  assign axi4buf_6_auto_in_ar_bits_size = S00_AXI_arsize; // @[AXI4Compat.scala 117:23 Nodes.scala 1212:84]
  assign axi4buf_6_auto_in_ar_bits_burst = S00_AXI_arburst; // @[AXI4Compat.scala 115:24 Nodes.scala 1212:84]
  assign axi4buf_6_auto_in_r_ready = S00_AXI_rready; // @[AXI4Compat.scala 107:18 Nodes.scala 1212:84]
  assign axi4buf_6_auto_out_aw_ready = cmd_resp_axilhub_auto_in_aw_ready; // @[LazyModule.scala 353:16]
  assign axi4buf_6_auto_out_w_ready = cmd_resp_axilhub_auto_in_w_ready; // @[LazyModule.scala 353:16]
  assign axi4buf_6_auto_out_b_valid = cmd_resp_axilhub_auto_in_b_valid; // @[LazyModule.scala 353:16]
  assign axi4buf_6_auto_out_b_bits_id = cmd_resp_axilhub_auto_in_b_bits_id; // @[LazyModule.scala 353:16]
  assign axi4buf_6_auto_out_b_bits_resp = cmd_resp_axilhub_auto_in_b_bits_resp; // @[LazyModule.scala 353:16]
  assign axi4buf_6_auto_out_ar_ready = cmd_resp_axilhub_auto_in_ar_ready; // @[LazyModule.scala 353:16]
  assign axi4buf_6_auto_out_r_valid = cmd_resp_axilhub_auto_in_r_valid; // @[LazyModule.scala 353:16]
  assign axi4buf_6_auto_out_r_bits_id = cmd_resp_axilhub_auto_in_r_bits_id; // @[LazyModule.scala 353:16]
  assign axi4buf_6_auto_out_r_bits_data = cmd_resp_axilhub_auto_in_r_bits_data; // @[LazyModule.scala 353:16]
  assign axi4buf_6_auto_out_r_bits_resp = cmd_resp_axilhub_auto_in_r_bits_resp; // @[LazyModule.scala 353:16]
  assign axi4buf_6_auto_out_r_bits_last = cmd_resp_axilhub_auto_in_r_bits_last; // @[LazyModule.scala 353:16]
  always @(posedge clock) begin
    if (reset) begin // @[ComposerTop.scala 171:22]
      arCnt <= 64'h0; // @[ComposerTop.scala 171:22]
    end else if (_T) begin // @[ComposerTop.scala 178:19]
      arCnt <= _arCnt_T_1; // @[ComposerTop.scala 179:11]
    end
    if (reset) begin // @[ComposerTop.scala 172:22]
      awCnt <= 64'h0; // @[ComposerTop.scala 172:22]
    end else if (_T_1) begin // @[ComposerTop.scala 181:19]
      awCnt <= _awCnt_T_1; // @[ComposerTop.scala 182:11]
    end
    if (reset) begin // @[ComposerTop.scala 173:21]
      rCnt <= 64'h0; // @[ComposerTop.scala 173:21]
    end else if (_T_2) begin // @[ComposerTop.scala 184:18]
      rCnt <= _rCnt_T_1; // @[ComposerTop.scala 185:10]
    end
    if (reset) begin // @[ComposerTop.scala 174:21]
      wCnt <= 64'h0; // @[ComposerTop.scala 174:21]
    end else if (_T_3) begin // @[ComposerTop.scala 187:18]
      wCnt <= _wCnt_T_1; // @[ComposerTop.scala 188:10]
    end
    if (reset) begin // @[ComposerTop.scala 175:21]
      bCnt <= 64'h0; // @[ComposerTop.scala 175:21]
    end else if (_T_4) begin // @[ComposerTop.scala 190:18]
      bCnt <= _bCnt_T_1; // @[ComposerTop.scala 191:10]
    end
    if (reset) begin // @[ComposerTop.scala 194:22]
      rWait <= 64'h0; // @[ComposerTop.scala 194:22]
    end else if (q_r_ready & ~M00_AXI_rvalid) begin // @[ComposerTop.scala 196:33]
      rWait <= _rWait_T_1; // @[ComposerTop.scala 197:11]
    end
    if (reset) begin // @[ComposerTop.scala 195:22]
      bWait <= 64'h0; // @[ComposerTop.scala 195:22]
    end else if (q_b_ready & ~M00_AXI_bvalid) begin // @[ComposerTop.scala 200:33]
      bWait <= _bWait_T_1; // @[ComposerTop.scala 201:11]
    end
  end
endmodule
